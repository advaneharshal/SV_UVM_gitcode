�Ii2�*�� É"�t�d�EX"����,ɖr�<66�%&ET���0� ~ Y ����EG+l͍����U���1����#��d����{H���n�g�<��n	K������c�xSq�ݾ�<~!|F�Fҡ��gn nJ����ĉ�1FĀ2�EJE3����ddɞ��#Y�Y���]W_�nAj(�B�u��CY��������|�I��O�{x�@���sx���p��jb\�P�qz](���z����u���87A̗�h[��MU���N�)<Z4`�nct�g;*�
�f�W��O��`c���j��]�T�+$F�7�k�p��.'۔�B������Q��`p.�W� ����@��ed4hX���aو�P\X�œ��"O�%C�����%hO���o`�>
p��z"@/��?��� Ss}�p���M
ONO!�f�w!~l+�fko�?�_{F�9�{��$6ٚ�������:v'�Pp>���;�윙U����c/P;M�����[���A:: �e�cbx05����kr��~�\�c�+%�/���1%@~ȭ����t7�@�|b�L�=՗��^:�&��"�7�υ(�/X���-�`;���oh�;8�����2/�����4�$��}��j�X,�~T�O����(����؞w�˻s��[~���Zn�*Sr�Ք��}�(J�j���h�֠ط�C�O��1�sl�H]^t���3��⡞�� ���Id�Uu��~��I�� ��y�\Hm-O�Rt"C`+�����G1����n��H�
�H��Vh�^�m><*�*���&W���1�Ȁn��X�����-s\S�j0�9����4t���>��!�d>W^3�b�_'y�ڕ�!roT�\q�'A�e)�۸{�.�u��(w���S7�.�,%���+���>g�\�կ��J`�ǌ̓y�
6�p��^H;G�+���I���ʡ�k�%�0�UG~Gz(6q*%�-���ZF����˷=l;�P`��Tܛ�����s)b{�y���p�)�b�T�֩ ���s���H�����<Vt���%��t��=&E�YEf2�xs�&�A���CX^�g0K�mrEANiV���'��ܲ��2�5rͫ$!�S1���	�x���6��g�y��^��%�J-{�2Z�
���sX���u�ň�wf���k/�05@�~��}O+��`���(�!䚉�v����v\ñ�|�����l
���@����V���a���c|�@��������N��~��P���+T+�u鋨׫�1s����}r��!��7��
	Y,YGidx����\LXQE����#<�[�ُ��[ﺈ�&�zk���L��
u(�f�$!���6	�)���E��6�*M��.&3��UŠ��J�:G^L���M˞�Q�:%��X�Z^G(PGƞo�,
�
�j"�}�ÏȂ8B� ����B
��Ԝ�/�S)t����t%W}W�{¿��-�����|X��d�o���fZ�V��S���b�����x#�c�/n�����:��?�����a�s�����H�OLz��l� ]���8������S/E¶~��b�I���w:��zm}�e�<e�sp0$�l���ϝ�WO4�}��.h�?K���#R\7�3��BL)�޷ܯQ���Ven
�;ch)#�f�������||/P��/��>��M]�!�&�.�x��ZnV�y���։�F=t��No�B#�]QD�qo������&��O����3�5���JéM��씇��7��E�:
n@����¿c��Ƣ��&�l�,�[Nj�FG�u���-b�཯	�(���A�Pk~L����=o��3L7u�"�~��`�3��>��T�ֶ�������g��r���#GN��zo��p��\�^�bf�X��'-�Ȥ��3> �iXb���MDA����R��k�C�U����������a\���x�����UI�r���gX(�G�L�ʳ��n���g294bu���Q�G
c{;mr'���8��S@�ە�}t���d5�����z !�+Պ�р?9\�,J-:'����)DY�{�P�.�2z���u��-����^��yo'.7�|�s�_<�=�iW"u'Mp��h��^8�d^,���oI+��ń(��w�as���)��#ry��NW�^"�עQ���̾�H�,yc��b4��D���+D#��i�x�M�l����#��M/8f!�ȹE5�v�'��I���&V�|>��X(��<��u����ܐ/���F�h��gN:Bx/oF�B�s���RL�J
��W�6��Ǭ��p�E-�|��j�5�=Q��!a���]�j�����^}�7���<����p��E8���r%�KXKMn�L؞r��Kyb[�Y*R�i=me>̀��Tm�ꯠuf8]u��Z�m�W��^�OC�K2�[�:��nIsA�j8�2x��:Y�5�g�8����ѸNH��yW�oE�x�� �w���d?�	E��$qQ!U��S\�<I���Rt4M�*|�!�A��Wi0ʽ7CL�L�댭�s�i�-�(�Hrt ��*�r�{��"4.�����.��zy��Q�(����P��aPB�w�r|�����z�G�����O#sx_P���V�a��{��U���#������Alk�)��HѤTiÁ� 5�LXu_z4�"��Qu8�"9���LRW��[����c�Q��F|�{Q��ԺC�%���+������r����d)�@����j������-�A5���|�:��:(����8���q<�1G��M'�)�Kv��$�
N֤����ͻ�p=ݭ>Ua��"�t�Z�BV:+��P��j/��i�wc�4���ɱ����t��X��A�,�'�+z��-|͹�������Ӕk�B�՜�.u��'4r��4\�~�o���s���7j�o��&��Z�\�M�����1˅U֖�t1�.�)�b����!)�B]�.r����rĩ�f`�q%b/k�ީ�#�L�ϙ�mN_�T1��U���.��H$����>@*�-�]�N�f�tP����K�Wt�Y�pMq!`����� s�&!�`��b���N}Sh�#�m�mn�16�Q�vS��>�w��Ɖ���4��ﲾ�ks��=����)@c�P�D�w�r��G1��%�U���J47C�ژ`�|��I	���3�&;l�׽�3ԙd�
��%=�38C~Ȅ��E>34'�`���q��p/l�Q��G3�� �=����
I��qj��P�?��_VZ�k�ܸ	}�GSoA�Pb��z֌l5���������YH0�(R���G� ]����r��!wè��t��&������(n�!�ՠz5�>] �.��l��R��[Gp��18�6X!u>u��v�t �[9.(({3w�S�M�E�/��Ȣ�W��mz♐��S�Z�z��9��֢R��~v����=��M��\��RۣCᗫ�8\d�5�K����{�7R���;���xa�vm�)��=p������D�A4����pM�x�%Q'�Z��~�F2�),Bu<����0�����jQ7f6?/�$��$��O���<h��<��Ůd�fb�I��h�n�� ;*x����jw���ݪ"�E��7N��p�|P�mҒ:>@ K��Y�����H� W�*CaW6H��r�U�Ǳ����n���n���G���y,~�p�j·�ڔ�2�x��!�p�׮b�����8j;�
�1��V�鼼�W���N6aw���i���S�x��a��ޭ����_�2
� ������p�<��R]�,��:���D�H	��鬿'�c�ԡB�.��e�
x�Ri��֝*8�`L��GK���e%HOOG�6����*�[�&$K���5Ξl�L����F�4��M�+@C��6�A���F��ʇ�x�L��Y!�<�4]$�X��-��.<�	��|⸦��]�;�.�"S��@H�N��F�NM���&ʁ˩\�w^�e���%W)/`� 2@�k�] �4T�G5Ÿd��� XY��<�!	8p�~!W�MZ~�֭7�zR�3V�* �����~���H[�����M��Y����|5b,ㅱ��[>M�=��D�:��)��e��%�������Q���n�+�A�љ_�X��C�ٷ��X�PY��0^/�X�Ywklъ�]��z"�����rR�<�Otc���� y�=�q�l�A���d­�Hp���O,P_)��Og��Ǉ�=v�S��!�q#�M��-�cp�	N�#������V��\`�~7F(V��H߬�x��ZrӚ���� nĠ��?�����Ow��1^�E��������K~-�w�V/}k�p���� ��aVb�@4	�~�Q$%����n��(�k���"'�K������p��7�	*5���C�|��(��lhZ����v��Vl�KO��B��<~�.ĳ��xN̂r����hzS`W.�k� M̌�+���2���*�U�f��g��ct�Ty��#M�XY�ڏ5����$;�0(ls�M(��i��n׳`�ىs��Cڜ��P��I<�����l��<[�`i��D���z{����&�E����������(�/��(ү-��(�;���O6ux��;���p��2�=�Qݐ��d�kI�d�ھ�����pV���,s8Mz��0�B��PX�_���-�%��J�'RZ�9]T�=G��6��q[eeu/͈e���V�K�Y�"�>����"�	yܴ��m�s���+�gc}�!�죠��2 �_����\Р]a��/]έ�"�Wh�JCXM6�w�b'Ce�ZV�K[M��;����}�Q�}�ٰ!W�N+%�H��5�J��w6Q��)��D�f(���09FixG+�VG�a�n1f�Q��͙�t�	β���ʬ)��̢�������h���	�Y��p�:t�f�k[F-��X�jO��'��yˬ��+�yӶ��ceh�#o��A9��	oi��],=�ZwSo����^$xO���U;�4GC���v�7�42������ń}!A��D�ݓ�J�!�y`5�������+Q�e;���=v������Ь���Y�'QL19
��ɉ�p8�.*4
abx�ci������R�Mc�1��Z�[��zq7#��N�f����?j�L�b�Ǻ��y�A8�ݨ쒝2��_�N�O���-��!'*B[���W�\�-�H�		�M�'4��T	?N��q�I���m)�f�ͼ%�vn���i$�{����k8j�M�{����4�ܽ�� �_O	y��fh��t�
����6ki��bUN�[	���v��~k�땍#zs����<���KB�^���I&��ʥM�fD�
��3n[���-o��d/S���*�.� ��܌�M�֧7�*�D�Ȕ���8�]���HCخE��^�
�߲}��]�e�&�H��^kO`:�ʴڄ>��Rt��_|g�J+��A!茻d��YW	<��hѬ�!�R�8hN��g��2�"w�w���|��E��St�Yj~�������`En�����B(VVQ��0�I;�Nˁ ��h�IHu��~�?��ye5ՆF ���sw��طR�*� �q�K�7&+ ��Ə_U�j�-��1	���Q������+|װ�h���b�7@t�K���>�M����s�2���q5��I{s�@��z�βg�x����ҏ�o�L�c�ރkw�x�#�HS�Y��|w�&ͭ?�XJ}�a�mR�~�fm]�XxЙ�I4<��n궷Gx������c�ki�h��02�_����ע�FO�X8�����GQ�y�|�'�:�M��v�>���邃���}��7l�(.�T�X�2����W)�//�m����C�T���-�A!`繆tYG��f@(H�)���7\��Ohs�I�Y@W��bY\�Bsǔ�rh:����3Ln�Ӫ�^�9���gǔmJ̒B�	4�;U���q�.R﮵j��y[3������Y�&QqL�1�S�tzl��
���bsf��5���n�0��u#���FRG0c�t��pu��r5���P'c�C�y{�O�>җK�.G�F��w�������oJ���1��`����0��uqp��ZR+<�sw�ۜz��j4��i-fր+@, �t�k�������h/i���V�w^~ �C�
c����L��s�<�C?=>��X�� J�t� �u�)���"����'.�j~shK��^�~5�����i����X��$eR����v�v�����M�{��K(�h��)I���}�K����<㔡��dJ���$�J{� Z��RN]�k����UM�1@NN��^�B�8���q���)�4G�����2�rv��.J9P����/1���v/t1�x1O5=DP�k�%\ч�
^������ll�e����s���Á�I[��3����]	S�`��"?�U�{
��T�!c`ǝ��~f5&}7.����$S��5���/i�w.��¬�Kİ���ZaL��F�"=�|�P%��"˿!O��$Ȑ��	J����?��uE��<� Z���c&��c'�7�>�&f?
Z
�}<D/{hU�۴�`,OQrB=��Vr�pG�R3��60tݐ����Sw�N1鸣�3~�{M��o�S�O���5����M,d;��>��j�)3�헎��� �.W�J�~r��]"�2�k|6�O�P�=����7��8�$��wI3
N�v�k��m���PMWz��"L���Q��-�z[,L5�=]���'�����̬���y[Ay]ˋu�<]h"��4 �*��Q����M�`�$�1�HFm����&��Fo����]�¥3r��^�� ���^5��à�o�Ԑ>��c�Qd�TcC�����b��o����z?��`�������·���Jᦎj�@�z�-��6�+�ϑ�ȃ^788���4�أ9���RK��[�ĐOF��q����$6�HK2�A�$���hԙGHy�

HiC�i�u�/��A�S�xەsm� �S\�C�U�]��n�zR���y�ܚ���&��'�@4.}t[2??�[#���jo�@��K�S��b�t�q�:�����K��R b�����iZW&c�b| ԯ��A�롴y�u(�����/������\�1+DdߏsN/λ��
��JH�2�������D����ƾm�qH��um״��UW2������q1�rt�R��Y,,��zel�??;��9�l�SU?oL�y�+��]/��Y�S��R�L&�	K/xwp�����7�抇31�>�0E�*�Z�@Zer�GZ29�0������DZ�ݍ�ˌ�;�v��a�#�:���=��х���pѭ��fc[��h���&5x^�2v��*Ξ3���?ӳ8l29��'�.ɉ��S�8jr�.B� y��'j�$3�^ڗ=5�������'T33���6�����g6���t
$~�I����I�^��"�e������E���@5tN���Śé�#C	�f��a�Z���ۢs���|��'��O]S���/�i��t%��A��c1�&�t�y�r���9ΕT�|L�V�b�O��79���uiR:e|�w�p)�]�` ��Z�2�?�8�8��j0���rw*OQ�>���+Ì���]��C�o� 8z���V�������)˒����r�a\h��?���q�sO0ߍ�#4�9ּ�e�y���B�������l,5�ON�>񞝲�J�u��#�I����T{7F�/1y��?�Χ��'�=m-�t�P������/�f}�,��ü�Z���	��-t��k�lU�k��o�hkE�l?6}@Z������ �(G^ĵ�%x^x{�����+|����u��t�I6��b�Ⱥ�Di�����ɐ�)��8��D�+S,��5-QЋ��$����2���AT�z���ӗ�d�e��9@pdl	5��[8NrͅA��x��3�w��4l���8��=��¼�T��Xӧ�P��Eٍ&^(&�Y?L��{��5Pj{�
`���CjE�４�Eq�����U��=b��(�� RDɝ^x� ���N빓ӫ �_�<пL�>�g�Vd��f�ʈ�����I0(�QJЉ�`��}m��k��o����B�Uz��;���30�v�� )��'$7��e,_L<I�zM�'���\�=+|4s�$�.���=�V���SAI���tﭏ|����#�߄��
✕j����xB�*��:�}ek���0 ���}iH2���"��RiJ�0i�X"�[��6t�D^�]iAP~J%S�:s��Ud י��q� Q�����}1Q(&1��7�#c�7��0��� ���RIh\`�>���ġqu�r�Ɯ�SYin�� nu���7�y��W����gU5 �84x���3�l�N���?�:��v�\z�?�$uGJ��}9��/'(�����H/������S�7<s:�_g� B��2�=�:����@>�]�#�_�Z[<M��c}˪�������g�r�̌O���01��b���h(���HM@^lY����Ǉ�_D�~��t��̡��Q���d՗�S}B��9���).�uYj��h��޶��vt[LP�ɦkV�.#��Oy��*�����7�`�I�{kզ�!o�VcPR����L�u����m�N6�O_�ꉚ�iڜ�F�m���`n�/�*���S/��e���O��o��6����}�9C���6�r�
k���=�����%���P�������U�<�>I�O�Gg`S��HB(@ YEZ��2��?6\�k.����!�1Re'")m���!�$�A�1���Z������C����z��
�qPt���0��`�Q�o�;��0+gq|�J4���x)�YtxO]�Otr˄üX��y9QZ:*�^&�W���.�O����?\`}�P3X�,��w{�����t��������ǫ�P>��������R/��y\gE�|��b�,;�'�6���b?�jc���-<�v4���R��S*z�=v�Q�]��.��/�#S2��^�
0����cx����F��7���h�am�������m��Y>g�m��N�d*(6-[�_"I]q�O��Q���p;����4�O+v?&��l!�#sj,�
����xK��C�$
|����7��� �B��4a��zS�ֹ�y@3��l��w�]�{��;�{��M̦��8(���ɼ���e:E�w���2!q��b�����ِ�$�`��D�����N�j��t��R�օ�"�wT������pjݣ�R��G�E���z�V���_o��Ű*�7���)�Z�4'��Z���dV�w�d5+�;J����0&�������x7
x4��"�i��YJ�%?����'+�N�Wҕ`��>�F5?���<_P���6��������M/ѹ,�9�g��fL8[����8]m�@.r�ȶ�4p�U�?H#A��d��;�z Ĉꎝ��gQ~���+< �ۺ���$^h� ���n�5�Vq�����2$�t�Sp}�`=nʖ��F&}�"K$%rȄ�9)�����H�
� ���h������&���1	���Q�t��<� אqrO(�R�'~l�I�.iQ�j�(IG|<1��h��BuQ����3g&�?w�~V3�?��uL)(P��SWV<��CWAFa��`CF�{֩j�'�]�^4F�d���I�@"�:0�j�7�Z�����ۙL�4���E7���!Y�?Y�O�^Lx?��,g:��|���\������:�瑑?����Ff��cl�v�_$���}&ӥ�il^ۛ���S5u���J� �q�6h�`u��ϤY%��\�����R�g�� ���6ȂKȒ/o�FJV��[����T�	;P��Tn5l,2(�@kO�T��A�~7��R
؀��\����S�l��՗�����*��2vmǝ�;:��H,�m�~9c�_�w�L��)��v�I����/�g��,�1�K��~�꥙��X��0��#A-�?�*z����_�/�W쾏�e<AlP��b��Ќ�n����WW��f���b�,bd���*���&7����[�u�1(mm-�oE�g܁�`U�.z�`3� �B�_�F>�	�i���Mg��G������85�VwR$�B.�.�
���BZ���r�H�|���VUݯ��X@���L�M9V��f�����硄~�{��8�7�*��V�bt�si6ҫ֨+#
�55�>~�ǻ��:�d�~4�]�%KA� ��2�l�>��3��r
�i��s=Fʝ�ﭢ��9�_,j8���c&y����'`Po�f�h*�-�r��LuS3��񚽀Έ<��)�LX�������P)���2l8K�z���'"\[(��8	����ٷj�|�!�CXD �k���sʻ�v�K�qT�h�XE7H�T&/��n]c��@��L��ו���� l�$O���V�5������~t.>z�-��FP��[����)�ՐK���WEb}bu�[��jg��[������|��hܽ�t���*�4���MQÐc��}G������7u�k!�q+e���]T��K��շŻ-�I|� 9��ƺ_'�FL�Z�*4�B�K�I4&���,X#�[�-�4�M��R!B�ՈVv.�q<���_W��Қ.�Eu_�V@��������*|���h�OZ�t$��v6V�|����~�deL��c�(E�3<ɟ�"�($�F#jI�h���M�Q�nqAJ�x��#U�Ƕ�4}}����yt4�fUy����>p�r��2�ǎKi����Ă5��f7<�=o�6h4I���Ƅ�[$H�okV`�*��K���7)�Bp�(|�AO�4b��tԧc.z��AN�E$_8�3�&�����*G�����%Ք�0��8�tӹXr�%>*����X�]~��Iu��@i1[p1�r��M�%�[��'q��ȧ&̐e$aT],�?�=�20�ɔ_AH��܍A�{�Pm������	��4��;R5��L�^I������D`Ϧ�3�r�x���� �n��QH]m:��E����O�R�`˂�jx	��Bv�����| >���[?���*u�o(h���}rZ9Q���X��1B��#�v[�u2P���ۂ'��8"\v�Du-�AQc<�K�����ݿ�&5�;�W�=��������R����s�As؛��BRA�GS�s,����ї3�����
�q��5MfS����}i��zȕwS��řJ���%�:1r9�>����ϥc�s�� ~�pQ[���*+�S�l5�Ô���r��H�?pNO�S��+7��ARD6ZY�l���n]͆�H^�%�@~Y�#M#�ii�9/� �Y+���ޠUiŻzE��V&�H���r�2auXo��e�p�ةM����YX���1#'2�t��-��i� Ǽ�P>">�`�T�55�,��Q�^��_�?�,�����z��m��zۉl�����7{qy��>��q�4���Hum�f;�,�5�Lb��L\z��+2��yѱ�uЙ.6S+xeE�+�V�A�,��@��=`(|��n��L�l��P?��OO(���?x����X�a�~���}&��i@�7�T��k�:�ԁ�ح�:�'��c�r�%v��Y�Q%�`w"o���"����
��9M秫��Ʃ\�޷:��uǡ��;�t�B��-SyQ�+�J�ٌ*2��ݢ�H���,4�������~K^�l�SO�)u��?Z�I�S�CpQ�+�(AՏŊ�LS��O�>������<�.Yu���'GT�m�����n
���lᐦ�LN�����]�K@V8AW��m�
�$B��R�T<D�i5�G�Z,u����)	��G%�GC�3���a��a��/�"\�A��D��b3s�Wm�oZ�v�Z>ٴw%������yxnv��j�h�7c`�C�ynvj��v+��vR�#�:��e�&sޚ��*͟<~��"]`W�	f��J.���Iκh�m�S��U����y^�]��)�R��j�.�a�,UC����7r�՞�V֙me$��D<3��{� ��U��X���g�>�ϐ���2֧���9��t�B`c�K����a����Z�h�Q��݅%}g4�+�`.� Y�{��E�g�y��`�B,� �V��8
����(^���� �H��IŐ�v��-�a�"c-ӝ0�0�"��$��ָe3v�L
�@��P�{|�I��� �*E ��0�6�-�bQ��X�Tc��coΎ9�c��S�~�=�hп�n�y�jm�nbQa�e��c;���	ӽjm5r�Ka��L|���Pv2P7���c������#`t��5����%5m�E��BU�9)!:��iR�����ܠ �]pу�4e��X���k{y�#X(/>��޹���xГW�	���
��M����-v�6eީ�ا������պiV5VC�� �[�T8ר� �=e�Sw�J��"yY��Cֽ|K���Y�F8�H*�Z3����F�'~|9�:p��^rX��+��:��F*C`v�z�>���8�.� $���%�6���r�<2q���x���S���.�9��M�X����b�2���ll�,�o�P(�?æb����'�� �-�P��������bZ�akX���M�5&�t�k��~�e )��N���	��k���~��a,"�E9*������#�ﱱbzQk��(>���K��w�(=<	��1��.Gm����4ڱ����0dh9JRIŶ�%�4hƗ8��$U��dS�ݶ��)=���3ء[��^7t�$���ρU�%�ʘ`..�t�@���o�Z�z�]�^�ɒe��rV���ٝ���X���T�7:��#�j.�����Fc� ��elc�V��.(+���%�7��7��题�����o��0��-xe19��3*�6�<�;9>�i��a���O���i�KPD�j���	�16p�S�b�50�Δ���cP�j�� �̅��DuN�!2��c,�,FzX �J��21C�>?�^w����f�W�SLh2 ��jN�EP��ꗃ��G�u������H�K���F���~7�u*��_�*>47H��*�����U���/�7��I��tĈ������cXlam�����9#�^�6W5nFd��>!X�?�1J����M;.��y�	wd���+�XZ�DB�x��t]�6�&\����1�Y�h�r��FeL}:�Սؿ-׻,�b��.j*53�%������
D+�H���,�U0�V(}�JpL��?v�5]O�?�K���s�6�������k|�<1�m.2(O�XǸR��O�R$uf7�e0�\Y>�r�)�c�7N�o.�.���4�/�N��h�D*�j�]�9�Iw,��67����5��)��_���u�C������1;Lx���}^���O@;4��
-]/u��`ߝ����h��:�`��I�N�.����z0�wZ�h�[3K�_Yb-~B;@�|[g��,>S���hΣuT�n��[1�4�oq��%�c ���"���>�箅�0fo��s�x$um��������o0�uU�'��JN]�G>�e�0S�9��%����x�v�|9�iQ3�ܮ@hĿ�V��ޚ�lt���J��ASS�_��#��������w��oژ�U����&9z;-�V�m�3LN_�0�uu��бJ�	ұ��1.X)�8������c$C@On�	հ��2�I� c�5��k�oVI�j47L-]��h�H�X�W�����yнaO�D,�� S���	9R�w�C��Μm!N���C�px!�ݍN��E
�Љ�%=ʼ�s�U��+�9��ߞ��r�7�p�ޣ_ԦQ���t�޾d���k3O�����	k��P��]l��5b�.k��m�G��q_��7SB��C�S,ǸY�m@�}��y�7�e��L�fƾ����ÿ���j8�,9~���Q�����(��"2�F�uR��
?��!��� �L�<��(`�
>\��`��;b1#�t��7�6R&�iX~�ձժ�D�i^��Rp��<É�Z���	yL�:$R�r�0��t�&�A�	���@������JJ�X�9d$��p"9�����C�:A�p��]���U`<K{dt�a�\#8�W�X��IB*H��{��~�*$�$�:oH���ɵB?TR�Ê|�x���w_6��6��Y�r&W�� ��%�JA���U�9v^5iM�T<�)��9�	�����Sp�����TҨ��90��N*�,�������u���q����}��k��1�S}ZFο[I���M%�+θJֻT�g����*��������'�kϞ�a�S"��K��b2���m�9��-����WP�U>�x��i��\!>��V��+�R[��I5�NF12(�Ú����E�-�f�����Ԇ a�`���b���ơ@����U��Ф���V��V〷��9OL/#��vg�	��L�|�\@χ��M�;�G�^օl}�SV���e�[|FJ�������.<*t��*`OUSm=Z�dR+$k�$� �vr
	�D�x���D�1ұ��YZ�ݘ@YBG���˱ O��^?ջ��������O�K?-٦���u��)�\̘Occe��e��vB-lqOZh��y�㙀5V��̚�N@T�Zc�ǒP�d�p�	y>���6��Dݍ� �a'�`9ZE�D�hv\���!ڣ�;�:o��w��R-���3�ʕX3��❚ ����[	���H�@��ç�����L��ȸ�w-�_1>5a<o�;�F�d���I�%��')q8 ��d���t��g��
�6�ciRh�����ْ�)P�r��J��\f��t�8L]�����r2yi%�+À�y	�h�F�<�p�z�H�}(#܋�/��:���}�#�$�a�Y|��1+�6��#��Á��U����æ�L��;cky~��x���%qR������B�qf���S�?ɂ�Zv���g����ɵ˱Qi;��^�׹w��]	���Pر����JE�x1���Z�C�Y=��"H�B�E�J{|�'�"�v��=;7�ͫ�6Q���i�f���ђ���$Ji��1�h��>m�8m��
L%#�3��y�ߙ�C��G2�N�6WC�̳����{ZQXa܆�~ E RC�
��tPz�3N�Vt:�|?�[�n!� �7;�-�7��!Ag�Kyг�G���T}�8?��u��N�,�7zf��������%x��t�1��� �b��ڝ��v��L�U��L�/f�k�F�d����K�1Q��N�*vws�>��Q����ֳM�3i�Тߕ���R�J��Y�1P�F�IT�.;Rۂĝ�z�h��GbE6s2b��	p�B�x�d�M�u�=��-��5�\j��-���_�^v ��3�O=/)�Cg�W$���$��]m|������A�ѐؓx���T�槑H#&>ʓo?O&TP��"vTˣۘ[P�,�И74n�Ӳ�fz�z/R���L5���G-��l{��Џ�p%�������![Ұ�a�f�O� '����ܧb�͒j�L��j~ΉQ����d�$?���wN�� b6�5�+)��\x=�`d�ާ�d�����þ�b.���Tl�3M��W���F�o��Z�zk&8�l���6�?������3����=�T$�������-/=6ɥ3���5Y���L�P���������j Q]�Z��;�O#5}���G����UGI���N�\�h��M�%�Q�l�a�ż��2��3��L�P�Ƙx܀v���5�Ҫ�$�\���C���{��{�������1L�x-�w���EZ%ք_�s�����	�Qc�2�<�n���&+���R�I�L�Eg�/�|T�?�Zm����*��[�l����J��ru
��1���/����G�N��I�1�-`#�s���m�%���ۧC�Ai�r&}5@`�!�	1��5���`���6gg����ܕQ�4i<H��\�$AR��nɟMK�l�&&� n�
pT�s�r��ÃH[��z� �A��.>ƛ߭-2��m<�EL�������9&q��a���Ȗ��`�Á�?^1;���B��w��%���i�H��R�u�8B@M�|t��q��9��Oh?�P#OϏ�ҕ�wE*xA��dZ���2�w�@����%v~�<	~7�F���
��
8$�Ra�B��%������!�\��i�PȦ��G�'kE�S�}�eF�}]����A�[�����.f`4�Xַ��(�",�e:|S�}ގ��������5�%�kVCI|�}Nm��㥓�1y�Cy"Bd�ʙ�ٛj�Vʩ[Yo�&�oȽ��$�+6��oDr��p=x�m��	�����hQm,��L^O�!���a�(|2���$[��ɜ�u�V��B��4s��!q��j�*��ǥE�֬��j�o>S��I�I������+r�}!�<�� >����j�~�_����+��΀�J����*�?Ya���Z��^���-��}�X�.��,��	&����#<�5��Ud�P��y�x��l���k>j(Xnў��}��YR��ܢ�mT�&�"沤����&�\����Ф�ዻz�:���:�0��
���p}����-�axNNW�Ӥ[r�pgE�Z�#[h4J[e�Bk�t�o~�����6Z9?��x�+ �v��O:0ˡ�HZ#L�uL�ؕ͒og1!��>Q6����������
�X�i�7� ς��R��8�u|6~���x7*�0�rK����k�����}�����~q�#
�{o�Yi�m��}+/��k{�$�Vhp�X`V���/�fU���>+N���.�7}�=�J1ױ2xL�|I���.��Y$J�*�w�"�����	��W�à�,G�;d�خ���)�M�~"�B���Ȣ����3���j��m���H�O4#;^����u���n4��7���gn�F�p5��!�?C?u@Alor ���%�W����Jd'tz?�T%��u�qC.�����S�l��CN��kY�eZ��sւg��0��U�������_G/W���u����4��D�E�R�ws=�����RyCl[�x:�<� cc�5�dm!Nû��=5�XV;ݶu%�C��n'�������A�M-�'��3.�"��I`�}�H���G7���8���,�7�'Ԝ+�6J�������р|3p,o��Mb�5	(��7$���M�o�o駃k
�*�$�w�`�nbͳ������vk��{�b�<����_������
�
0�%�cS@k����m�kwL��Vl6���@D�@>�=�W�ڦv>�
�	���jٹ"�QE�(�(0�����(��� !w7t�� jf���Ʋ(��Ɖ��ү 0�'��d�]B�na ,'}�]P�q��jT��@�,�^�I����t�V�f�ߩ���9q�c~�U���wm�q�1�`��Lo�ŉcl�*mܫL� XO�<-�``Dt�  hU�ꗴ����G��Q����F�>*�N�S8�,H�|�|�&����J��4v4=as9�^r.X��\A��#O���?��D�[E��c���Z�ѕ�1�^��^0�Ȁ�T���5�\����VV+��<�G��}�:� �ʁ�{�P_��Jr�cS�>3�������蹛�0�CwV5J~b�M`��f��C��=8Ms�	�z��e2�Ũ�AVPY+���|�(v�.j���1QR�!$��>.��_�B7#�4b,�4p���D�EfJ��W�e�r���m��Zr���4�X�An�����o�+b(rd�O��X�݆��\l�*cji��{�*�D��0��ϗ���Q3�1=+�r��݁���9!����Ŋl�����c�����	�T�nR������[������.v�

O�\�X��e���M$�BMT9���P�<
99��$Li8zV&��\��H��t.�K�'��S
E�<�-��">�wm�j�sQ��!�.�l���:<������v|�`?q���r&����F1 AR4C�����26'7?�W���VDsC����{��÷���=J��b$���,aY��N9�O�P����j$=rƲ��$.8�˻��W�bY5�����o�Kl{P1�jE��f�G����38�
�ur�g�ɂ�i� 6�L⁗�^� ��-�1�t����꘮��Pd��558Ď��7lƭis� ��Ov�n�i|S�5$�C~���Z4�,��.B�<m�zؒ��G�t"#d�{
��(FIP�������Q$�m��bc���o��mp_sǀ���!�.��R��>�"A��׫c׿8��!k)G��=$�X��ru��d8[�5 ��v����<ƅ���Ӂ���=�}�ɨ��XP��"5��5���2 ��(M�<��~��u�&_� ,9d%A����H���o�'o�kryn�c� ���x��SVH8�	���XlI$�/���� I���l��R���8FH������׬��N1����ܩ��{d7��r��0������� �7���=�f�0#rH��N�c�(+�M���,E�#���]���-�*��Sc��é��r�O���8#�J���c۽�Kņ�ԍ�kxl���q�>�h�6�^�}�M�q��ޯ͊x�..���v�R5�4fT���6S�Š��Ć3S=s��if��|���(�g��H��32Lm�?��xo�ڌ��8��*�pE�+�'�a�;��x� ƨ���}�KoT��h9��l-�鄢�	�Zq0�P�?K��ƨ�W��w�s���n?|��Ͱ���Y<E&�?���SYy
�[��e�5�Ê�`;�qa��y2B���-�� Ki�k)L����������ʟ+޸J�mk�C���pqCa�h4��Zܒ2��=�b�qfs����}X@d2�T�^Z�,����tك,x��ܔ@��9@�M K��cQ�.�D�ߗG0�×߅�����|���M.0��-9�׿4�ZN%���^���`2r�K&e�^���t�mA��4߮j]��_�(�Kǿ!H)���f(ϒM�ߞ^s��F��%U�٠{��3`������j0d���$6�j*�t`���o�:I�Tt�ಬ��C���uw]�`8�M�z%���C�\Pq�C�������`������!���K��>��G~�Q�J�b-�0E#�����v�3��B�ȳ/��=uW�'��3�rG_��^����L8S�<T|��
PGds���s���`b��0�8r4�E�8��~��ُܽ�oǧzi�G"���0��9�+q��M�К�1�����L�(���7j+z���I�T�p*��.>��ܸ�W��@~�m٦,hu=��O�E�R�����λ<�-�
���v<�bkk�^�ڋC^v.I�X+a���m*K���p�I�ߕ"@1�-��j/���Y�$�w#��zbV_���f��'4d�*HC���?�~(���-�/��eg`Ԧ\�d��K�~��	xD��K�J[�ߪ�]��Q����X�C-"��0��e~��6U��n��{��h��<����p�OǢK��h����>�g!oQ���1�AS�����G�M�e��7D����;��s�0_��؍w/�Yp�FIfJ<�cY�"�T\�����q:�5(̸�45n�.�Mb�
�����p ��io��}D��P�$�������N���C��W���^i�C]K��O�~�0q��5űQ&z��~������K�����8��K�����<L�M�����?|�2�}�b�Ϲ��
�t��R���ȁ�<YV�0���i�
���M��2T?�g�~$t��g%sN,���pg��X;���n3;|W+�n�q���
�Ыv�%d� љ����n��J`/�.�4k�� ���1\�����:-i�ކ�a����b-i���e�3VwU�/��Wg����^�4�+:��ȉ��Ю��q�*ϴ�5�&��m���;�~���^LfSd�]x8�u9���=;+5�� j���K']G����/�	��{������#h�%:.ʄc	/wF��G��#E�G�އ�@��9r�;�Ǒ&�2���e{ߐ��T�%�!�E5{�zε����*_��H��A6*}d�4o:E�Y��OR��-���햓�4�0�2+����j|�t;�C��v�w�{��⃩��K���#���b���K�4O�J!aN1��q�+����
����U�IǢ�W�,8Q]��x��3��9,:r&I��ߔw�a�=�/�^�R���mє�^�fOVc�Z��D{���B�f�H����^2���~DKN�V@�����ե�$�k��>��91ֺ�_��/��:euB=q��HNn)��9��7s��GOYk8��m¯v��X�0b ��e���Ir8�o���^�����2�}����H���X�j�xƲ2M��
Bt^~*3$��٧k�s�3N����T�� B�Q��]6{�S;1 ���de�[����Qv�T��ˁK��ęb�"��I�~aDoۺ�Ax�
���� i��q�u"r��?~� sYK�7��ZsN9g�,�!0DȯY�[�%�_{�Yq�{�U9R�p��QǮ� �ۨ�I�u��<�M�1�O�mA+4���` jj<�:���7 =�Z�S/� ���+O�9�͆j>�W��`�+"��,��>�A�;�<Ǝ�ڜ��"qג�UI-:tCw�c�qx��E��~��j!�48l�'��F�ͨ���;�o�#�6�ĝY�JeC���u+��b�`L<W�2<�R0a$A-�KC�	Z�`�;X\䜮 ���l���}q����)CR>��x$�ROϘ7���F~�9��]�0F[ZS��f��������1��"ٖ&u��5_e5���5�i��5W��)3\=q|��+��d�ܛ��|�zo�uD����#�5�Y��;�^F0ƫ�*�^RN��Iޱ4l��f��7���MGү	q�A�	���݋f�_`�Pp�YH�a<�s�@��x�b�No����H���RXu�VqT��YA�Ң�QqFO��0#k{#R���aB����K�j����X����њ�`���F��'�@P8�*;F�[?8>�O�����z0]�L������jS{�ė��Ȓ�,��yy=�F�+���/A�����~(���D�T�fx�meC+Eco�)c��W,S��%��S��:V��R��
���J�T�!U�%<�'�o�k��Z8Ҫ��o�;-��qzhђPy�PƬ�d��2v��Ơz����������^�t>�=y�O�Х������A�q�6v��Oy��-�vy������`$ ���j鿩B#`ʃ����\t��ig�R�jz��u����<_�j����fgΤ�Y��KT�f&#�������{����#����3U���̷-Z��$t���	p��'�<�J��Z���r�����[�mc[:'ٛ@�ԋ�#�:�?z�ԏK�!;؆ Wq��x�o��9���̾�`�OW��p~=�.���E1�4�+����
e	S�Gt�rx�o�����6rW�h��HoC4s�.�1_MӖ��__����`��za��5#h	�ep�)S���<�^B;d�}��c*��D:	��ohb�*�� ��Q�ۑ��oE�����0&��֜C0�<p{rv��L���oR�<��$�#.� h�~�R��-�P��1��f����QQ����	g����-�g�c{{ZY��U3��k6K?�/�6��)��Y�'�Ahތ���L���,�m���p���AX���9LT�U��K��K5���5�H�������Ҏu����=���,�<�F�����W�S�>�\��Ayq��M#��9��1=��>�K��5�w��z�P�T� )Q-t���<�拐��U�E�ڡ ��h;���v�;G�@D�?X� ^�t���e/���n�_ާo.(�w�R.R�g�a���}��@��FėI��:Q+"��N	��E����x��<mN�<v!�rZ���d!. �yK��F��Fm�3��t�	+�H�X�U�i &hƬ�L���4�Tn�=
'��Wv�vL��iwà�%`��m�\D��mT�1a��@,�H!�7V��=żW*B��!��e�=��|Ɠ����hF+�k�Q�tZ��zmzv��ݕ�:���b\�=�K�uL�C`�'����>.̨rI�Y��5%@�U|7�	��Oj�T9���>�^�	H��$A��I4�$����5^�'�6[�Y����1�������}>�����%8�06G)��͑����������w
fY|ɒ�NoO��i �������J�f�-��Ķ�<��}��"k����'/s#r�{{4��w��`3�V#�[?������ ��%�l-��q��2r�w.^�t��qss~a^�9 �f
�.�	sU���AM2/���>���oT��-c=1{i�JD��!rh:^o� ^��)��)�F5���_�������vy�� ��w�*��{4�Ëb>�>��V����^y<|����A���`�2 1hC������G
�`ٯ�/@j�U�K��TM�D�i������g|Pz��ڬ�_���T�S��i�F�|@������J�avzB��%|Jڜ����	P~2�࢚{n���T��\�q���pu��ޒ��Q@	�����n���m��Z�S@Mَ�䚜��9�v��Hîte����u!5��諧��wmGxU��*�y �����oVTaKPg�jSq;C�0���f� ���uO�z+�
1Z-�Bs>0��d�٘�p��0���|օ�%����*�I`+ִ�`���t�JX�;��JE�-&��%74���ܮ�5�)+G�U�c��CT��o���ҥ�6�˹ù����L������0���D�Q�q�6�*��4Y(�(
���%�wb��8��}'�UZ7l�F��
�5��)J�e;��#ng����7P�x^�<d0�eg���l8��7ot�U���q
�D�kw���H�Y�1?BUÔ�Q��Ҕ#^(���������k�6�-	{��,�a_e¥�{� Ǻ���!��٭C5dk�.��|^�)�d�N�=�/H�T���N�����1˱
#%�Y.}�5]{��e�P�r�y��~Ρ�'�%�732
���MsG#��1�&K���a�������M�]�sR����ܒ6���9`�Dx���+~%�v�dK���ʳ�Lv.�3U�BxL�d�٬L%��51��=H�@E�p��Wq艊q*���Ն�?��V��w���)ۓNf�ı��M����1�n����)�#���B^c�9�*{��KJ�r#"�4��T��;~�aC�X�ؠv:��x�*��Ed�����p���UT �������V�aq�Ƥkįnn4��R�i�/'eY����?l�Ά{V�i��@��h*V.�ܐ �-�B��$�Ҕ}b������^�2.`�8�¬�uKo��sD��CA����Tf ��-+��u̚���!G�C��u�(���{�6�n�"mW���Ჿ�H�Yx��A������E��M��o�`�eu��[\"����%��F�(5��P{�Qf��{0�w��䤨X�j�i���.%��#��ݟ1�O��mV��t�ƽ������Q����l�z�[��OI�`��a&�Ŭ=�&C���cGB���d�G3.X���7k*�$���?���_e%��R_���lp�&k}�,�D��m��_=���"�k�OP���fhxG$�?�*�ό8
P��:U����_�"�A��75���d�*^W��MdF~:�_����9Ү4��p��੫��sy�y��Q�ξ���ͪ9���;����� �MeަaX�4��%�ɺ2w�c��ZB)F����c�5�,ֲ�f)�|���ƑEc���o	"��\kJ@i���,n�c�^[�D$�j�X�k��2�����·�V�(�KZ� y?�l�Eh���EԦ��շ�� R�8�9d5�d$�2CH@�k�C��{���h�5��9Y�L+�8���Cw�:����I���3�=���"!^[�����������IN�H�1h����t��fá*\31�D.6�=�k�{�p�k�p����Aؿ����g��%/-�y�5!�싫��2����ǖ�I7��ע�ûėvKc��Yj��ϹU��e��,�_����¨K3U��Lp��� ���zN��S"h�R��qw�[X{�p�"�I��l��HY��7l�-_�фs��!m+K&���'�EĎF�mL�7�y�<���M����)$)Js�	�b:����"+��
z�!7�L�t.Ɵ�p_�R9w�X�3�~�����G��}���|/�uW��r~���������A���m"��Z���2\�'��ۦ+23�6�}:��~�
���58�0�U�3(���*t;h�]���#�M@:%����| �xe���s>2R�� _ �b6���G0�RRY�ʛ'���ʆ�R.�C{�h���hiۗ?���b2�ai���dY>Δ���C���pr :I�HΉ/���ӗ�5�o�`&Xi�?A�[��uw�A\&W:{�n�!c��w_�4���\0Ǽ��$����5Di����µ���,M�R�Ƒ�{ԯ��M�[M��I}B|V��}�A.�`��A,��6s�>Q��\��y����8�;5��Bvb���n���.�����a�HngQ5U�*GoV�XI�Coj�|v��"���E�S��i�����j����c��Z^�F��MH�Dc�4�Xem5'B�/�QZ]�@0=^�0�o��\���#͆S��r蛐���.Fz��´H� E�0����bP�#����C��y���'�QR���\�t\F�Y	�<�S-#�܀��,C��/�9|�ra�lg /�y��78L��R��z��;~��f�� ��D{5ǥ��m�h�Tt��q$s��4�����|ܟWN\��u�C�~�K�;-�@��x} ƍ�?o��֐m��M���T��s�^�ϱ]�6�[@��A�X�-�[\{(�R=T�CF���T��K���W#}�J�3�`S����#B {�����`i2��'��!�T�I��N�|^�`�޶�}Ɏ%��>D�I�@s�˹���W' ,wxzt���	P�/�Ba��	x)�y���L������٨�`�z����1c���0.g_p\��S)PF=|p�O]c�{r��hySP����Q��X�,�7`gəf}2��V#��80`��|�^X�'��X2�h�x�n�Y3ǧ��Anm�ܮ:����&K�&���Xu�w��G��v�鼍�2���a�
����+3e�#C:K���LX�F�u�߇K|)�+&KT�Ǉ�^����j58"�i8����%��q�{������}������H6�{Q�^��6�v.Z�Ԓ�s�.\]C�0d����OP��\��?��r�6�8�s]��l7ї�l4��8��d�~��E��bGXt�0�)#�������@dZ��XEODۚ�P��h�6�, ���xҏ����� z?�E�0(ϋޖXDT}:(�a�Y��'y��/B���U�8;3��*���>�;t�狂3 rǤȫNc3���8��a��{s��
��tZ��=F��F�e��"�ǮD��L�����e�;Ef�o7��a��&v�v}Ab��D
�7��Ĕ��XDuP�g@���v������y�:6G��߀L�!0�"3Դ�,�YJ0� O��-���3%���J�u��OҐ�@����<<.{�{��7O��T[;Е^ш �	ܷ�a[�_�Qi��c�Ƕ�N���P�uog��7ޮ�-Y�y�6��y���v��i�{�veĂT���,U0i���;��'w�>/T����NC��d��:��g���J�����oam�}|�J2�g�3Ȱi���0�R��$��F�f���f��R!��o����"�[�6�u���3��l���U����&���,	Z����	��x �`fd��a�oe_Q���v����k���$�dT�w$���i0E�϶I����i�ܸ�����3����P<��l�{~/[����2�;ϕ54��_��WM�#4�
?[4ZlX��B-�c��B=��m)pկj?��#[�R���:Lk��
��j�`�&�~L�ڙ:ۄ��IF1��2��a7����~���R���ۺ{�Y	Ş���"Sh�N �`��!M+oܡ#M�M��u��t�ZS´^s T&�<m���W�H��'�]�S��Xz"��u��i����5�Qrs� �{�ƹ��@*�r���K<�ףÃ>?�_V�m��x��W��j�Qr�د͈"��w��{`���~SiӟГ� 44�OW�]qȵ��;}�Χ���"c��ͣ��$�&f�k�7���O��˶y41�7Q��Jy��=A�<����_Ɔ+��n��!����R���)����_2\%]Z��9��ƗB2�{�MKEy�SB�
	����H��|9e��vfR���N�,2K'���Or����F�nI��B`ぬ/,WG㣺U��6���"a��Gk���ɥI�,�ګ��afݖ��a���Ք;s��鼯~pU.~b��ꪰ����B,ζ������1�]	�w&J��ۊFYĩ0ce�VW�"�L�vm?Wo��Fk[w����^;�#�IN/��e�:�BBnJ*zִ��uH������k���>*�l`���!��K��P}�������6��y��������I�[l��[�� U%�#�1P��q�ܫ�#�g���7)q�Wh��S�S������Ά�/��Fd�/�	x�WŶ�4�pu9�P�KN v}��d5�Iޏ��|�N�x����9�?�wj5x�TD��yw�		IJG�KD
ad�N�����<;��S�s�ށ?Ǚԫ�����y���l\�g��#m����bc��[~!�&�����ֺI��O�������Q^W����ki�5�6��ouͅ��IXR�x�D�7]��)vǳ&�(M�����Ք��MS���\E;lL����!"��!*��JY5$������7��$#�U�i�p��p~�.â��Ԋ��4�/�.g��������1�c��_-����|N٠�;k��]�Q�X}R��9 c��(L����4tC�R�@k�����vD��Gہw�]�ѸQHR3U�̺�Oc�_'v���e��	�H��U!��b�VpgY���.�l���x���3�R�z̯퐅Up��H�*j�0�5�!�h��_E��������^�s��-��������Z6��~����lԍ~}��H�
�fD�BDZ�X�4猿 x�UJ�1�d��
a\���AF�%C�*�pX�o�)��-�S� �z!��Ku�C�隕�Sǜژ>������B�)Y�4��*3ii1b�3���ݾ+����R���� �hJ=������܁�Oq3�!�����ۃ�%�=Y�X�׎f{En�č{�b⏖EC���lͥ��*�`F螬�i}�E�;��lO2t��y�Ť5�T����S�?�0	�Ā���8���7����n8��2���p�֕�gw��p���> 	`�~l%)T��P�G�NHW��ϣ��St��&nfI�W<)�%{�v�����u�G0��crQ9³���a7�	ƶ��%�)����u�
�l:C�L�#V� � �5��ę4Z���G�zhB�]�K2���q�2��=��L�^k	�L�|ݥ�	��7Hr�H��.�\�X�ivx(���KL�t$���΅.*��}� ZMJ�KJ�C��޸=!�!A����t�*�W�n#n�@_Hz��X�ُqߪ�־t`�!�yDk0c�ݝ\hh�X;�n�L�6ʡrOt�<$vao�+�����Nd�](,UmU��ҫ�@���T{;	-�"%/���	69��k�Ʊ���.�a�������c�>l�B�)�� ����!����8��hQj�-�πyCc�V��:~�&���t�k
�G��g�	�֑xD�����b&�̦,����'+������r�@U/�<~n��F��&+��D}C�#��Z���±]\4y��6�{6��h>�1[}��D�j�tf�zE�\FDE�@ǈ�3��4��ߝ��qK�&�''\;��:��.wXi���^���Raṽyl�>X�a��l�����N��C'H�]e9�]�|��V/�g[n��߹�7��a�c��3�~h�+���/���߅�����wiO�"��,z���wȓ��_��׬��>5�����g<?Re�ߤ&TG.��|9GIq��aҽk��c({羞��QŢ�Y@�b��W�V^Z.C,�T�
���AI(�g�>L�噐1�R}b#(i�,Ԏ�xW��K>�i+ �g�	gv/���U~��&�׷A�����bq��w��q-�o�v�C%��$8&S�����^��}��j��)���K��b�M*���<o/�t�X�e�"���z|+�F�Y@Sy\%ߪ�m_��`��A��n�]�1���p���@�Q�ϼ�D�hmLGa9N	�+�˙��&��4B�x��J^����R��+�^�{��q����8kA6�3�}���`�~I�W!q9�Qfmi4�<���� \�c<�.�R�}\���)U3v�>�1^�*'FhWf�`�Y���
�.���mއ��3��;@3g���P��Spq.�� \P�U�ƤriE��iQ���4�TӒ�s*B�m�����~~�R�}^�y�/�7��]j������H���|u���(;����Jc�)Ș����N�cĹ������ہ�����.�PX�R��D�|a'"��a��d����G��*�n�`�X��79<
�+��N�	&��(~��@��/H@Y�!ӥl~Ӥvg�n���U�>�\@��D����H�7�����8���� �|�$�y��8}�o���^M�/�V:L�rΏ�5����q��.{f�CѨF+���}N�q�sn���F��E�H����!F��۳CP�V�7
��|�b��V���FxG�[l�'%k�Wi�_@,��Nh%�o�7�p w��ǳx?��E�C0���G��6U0�ӎ?�����WA;��ݕ`��#tkX;fð�j�"k��::c t�(����?�sz^��v�?�\\U������zZ�Rx��5��NL�֌��rm�N.@�Ե�:A���" Y�(�d������4�ce�O~����R7��/�	�rQ��m�X���@QR�P�u��-3�� rfE&�Q��H�����CG��Cx��:@�v�=�ӳ�@�{��X�t9�������?�/!�~�� �������vNyDl�<���L�>3��e��н�#�!{�쯹���T�ܟ����ӈW����,�LD-@�.t�:9(C:S���(�i,�ol��P�{�~T.�-�lYD��vs�����$��d�@`��K�Ѳo��G'O����)�^��|G��82��%�j�$]�#�b�����3)�p92���6�3��ƻ���=��5vd�	M9ۆ�fw�ɏG;u�~���rO����t^&���ҙB��8"��K�"߂)�ǂWQG��6ꉶ��}�����k`˔
�y�l'-O��+cQ��v��)�+�n��7�HO�3��`s?	qmw{�_wڐ����F_�_���a�����:-��<Vق6\��Ĕ~6`���Z����� :��x�>������}f��
����Q{V�<�_U�^��B�g���X�d�lgC8%�0�B��gq�ڸ��uf. ���j�P��n��q��j1D)�z�vG�W�����e3�ߒmͲ�a�[Zҩ���E���!��;@���#��	:�}
�R��x�wx���z��<��5�^������ͪ_\�+[Zq��
e}�B�ٮ�����3��V�M?�8�����-��j�=�=(��z�_5ʝ��,�
�'��m��N0UZQ:i ��s��;|���;�b����q��O�/U΃��E�<�@ב��s�
B�Z0z�f ��ZF`�I�ܲ��<V@ֱ{��'yp����f-���N5�L����k5s=�(�$�D�=U	7H����~��cx������ސ �gՙ\Ah�.z����&g"�J�ڼ��O�I'�n���7��l������a��^���O��l�%f���>�28��RQ9�uX��wH�Q���$�s��gg���qlk5���o_�k�9�:��e�`Y����fh`�&�U���?la��1�`�\7�d�W�!�����
��)��V���d����n��ix^��:�#��B�~6 E{�[P���e�7�[�Q�����DX=�;-�S=n�.]���Vs.(��*ƾy��?�u?����.�#�J�`��`@Q�$����\�n�]b#�Gb�0G��8n.i�n�K8�z(@4Sy���M��������7"r�Uȵ�u�z5�ز���u�n��mRp55�	��j�`PhP���=	Q�4�)�+�<��Vgt>g	2��Pm�Q,n���F��J󡚍���՟m&�=����M2�W*����o��c:�#�7��� �q�)7�{�b̡6�� ;/lp�w��+��F�N@��`�_> E��yd�ՙ��u4��o�h4�""��+�կ�6�'����n�N���=~>p�"�?̌�u{��@���4�D���7@��'E�ݛsy��4�5� 4ݝ<���4�������y�D��A�-����+�V�J�@���gL����TZb���m��4���t��wU�?���;X���/0�k�e
�hVŷ��1V'��!_�=��S/8�0UM�u�:��F	�5����M|����Л��@�N��*8�`/Raf����P_��k�JCD�%&A��˟J~d�R_�E6
:Լ�{�����w[9�<����s/���=U��g�M���s�la�]�#�T�X��:M��-���{}��8;��Ǥړ�/:������ZL�}m�%D._�4���>H{鳖���'������M�ִ*��v��v�2^+��N�'{Y���:�M����D��[n��X��� �;���}]B���z���<>����d=�zC熬��$������q�жD��7��(�p*q+�Do��|1O7�/���`��2k�Qu�������9p1嘼E+ɉ��<���k��+3T�@̃���'	%��u��$ǯ�#�1��+a�Yz���5b�/߰���U�,��ݒO��aF����q�x<e���X�S��L0M���\kG���1��x8��`��P��g��F)c�%��%��84ʡ�%��޻>���]��^$YNȼ�ؼ|1;��6{�v��W�L�ɞ��k�vP��n���x�͈nWᏊ@
�^ШAo�ny�4�1Ȼ��֓�L���j�����jAo���Ņ������.�����7#P���>L��"Ƈ7��O��Oԕq/���i#���n%L`T�!A���<��O���:�A}h�yO��1���U�,G�+����-�����Y1�|�~��� qrs>�r}��too� i�(�G�+�yb�u�6
Z�J�8m
�����1p��׶(S0�b)��G���R8�����]AQ��Yf��'��B�N!��fj��)��kE$��Uif}<uR�k�e�r	��<�?~�Ӏ�D�6T�q/T�m�Wd$H��f?���c&�+�
&�f֎�p{nN~���{�{A�+Y��x��5C�z�9�t[5��
�{���K����;��$\Iw��E�
�H�%��ݿ��>��Ǿz�>	o]LJ-HWd�a8����3�zE����6 ��h�f-����K_��8�8�`��4+��n�ֿ��X5R�9#N��}���� �-Z읙����jZ��kI��=x&`����_�뤇)�����4c�y�｝���[�E���;�����=n��ٞ����$$ρ]���t�/�/��,v��V�2ۇ_�oX8��Ԃ�(����V�E^�W-�)���<��,�B-K��� ��q�EP}�@;��A�o�J�v�	b-��y^�?�kG���>�ԷF��l���b#�>U
� d2�!�lm��}�� r�5��ܫY��%�_�:��`i�G�se�io�.dj���y���ď^E��Bg��2�D����g��F�Y#�A?�[�j�U�<�d9Ò¹�i�/�C���,� A]ˊ�%ޡr5��Cĸ,����YS������i*�;�����w�3�ٜ��a�ዏ�Xg�Y8������yQ%%;ϧ���n�� �D��wǎ��.�+��Dn���މ��M1R�I#��ި\��ծt�J�|]>�hM^��R��*fb��х�4���ĲT�`ݡ��7e�b�*=Ӥߟ�A���Oνv(P�CŒnR�� ����¦[���D�\k�S�̠�{���;-R �=$W������L���V��L���~�уSt ���n���"J�3�Z&���ڃ]x���QA;��[�X�#���ueK�e��q�NY�d��3��SҼk��t��>J�)� ��`�.]�x���^S���K߄d���7&��o��1Pb�[H�7�s��	�:����/mg��%3���'QT����^��.1u�殇դ���sGK�z��*�W�ݮ_��D�Ϯ�7��<b�	�h�p�QI�"�@9���G̅&�5+���<�LG��.c�/�H��Xv�iT�����i��ɩ����#�q�/Y$��mр����Gc,�J�A��3��Ʊ��}!�֚��.B���UKQ�b��{8���:�s�B.f]­K��Iz(G��O��!�����v�+�?��&ߪ�lUJ��qw`�$o"�ܘ�#��vp�4��nq���o{�����hWe��JU������A�8km��4\k�6����n&T�NF�캭)�6,Gl���D���op�2?Z�m��Ҟ�8�`���`������j;%͘t�<�A�����E�c�g�=�6T�pJG�ީD��
� �v��P,p9���.�E�%~��?��V�������������d��:C&EϩW���)?�C���S��}h>��-24?}��f_z�xF3�\�A���\��[��ſ�PПЮрZw��a��BN��R�á9m���ஓɐ���v�5Vi�9 y�����.��)���'��~ׅjz �Z9��t�Y�THZZ�SP#$H�E.�&
��%�g���e�����������y�l��k�dn�����KSn`$�AE�'��%Bz���J��ӥ�|27��bYH�h#�қ~���kOS7�a��qK��Q����u�)����_��e�՞����m�a��-a^T4#H�z"T�����7M[����g����\�Wק�J�PR��x-Y=����&���Q�n�!Ɲ2&�_�C9���a�x�N��d'�<_�*ЁΒۧ^R�8+C;�_�&��Ӷ0�Z2�r1}�[?)�̠	�=���w�JO�!�J[��2�/t��?�'����w�����y�R�ڇ�e;��j'��(U>���kk�9ϊ��5�݂�Y�U�X���n,���o�|Q'�Ȱ3e�����u5l�����]��.|j����1۶�e��OL��&� �x;��&�[׶�b.��LG�8��.�L9�t剚�>z�ݥGp�5�Ik�;���}mmΨc���n�f�#��Vz�hW��V�j�s�t�9K��	*x1�����hX9�:�W�c6^� d�^�}��
vu�fj�yg�y��b�$8�G��s	d��eo�vd%35��U�1�I�~S�vTTK�l���1z�(qx���㗹&H��Q"�㍿"'����u>'���y!w�vװ��>o@�������/P��:�q�Z�uO�z���͎l ����$n��!��5�MS���ڕ&�s��'P�������O���0�������y2R�����E]���D���D�B�1�dg٥������nNT�nM/�ʲ&���2Ni}mpGH�Ë_)񟖁�]^5!��뀥dʅ.��\擑��=+��P����}Y3����ee)H
K���^H `����c3��5��?\�7i=�짔���>,7�i�)kd8����#Yf�����0����H0�� t<�/�Fş��o��*H�gu7�M�����JgZqt�K��`?������H�}zO3�Y�Fn��Զ�J�����F��Έ�����{�)��*G�-�<���бJ�E*���^�JT?������E�Is>?� ˡ��a.Ŭ����4&�탵����(˻���Y�c���^f]a����g6��h���5ރ���@��" ;�S� �dy� ?~������htH6�LO)������j����=x.GK������c�?���ta��&f!�t x����$��`]�,}l��=���dĹ%����4��/�5�)t�
����I�>���v��R?C�K+�rvY�����L�-�uH�{�x{	��ׂ]o�(~J�\hI��$FNͤt$cE�?L���z�!M3�@w��#6������E.:�zm�B�eҬ���n�M�r.*�y6�x;�cT;3�ݗu�-����$Hy����ZMiذ�'�l�k�w��࣬ۼ��>�4e,5�\O�:�!Tck���+��Ez7(7klt����*8��R�$9Ziw�*��8��S}^��3�@�^��f�L��=�	��Տ)��븺�heJ�'ށ�B��I�] �%v��Ze�m��P�H�� ��'�|��&��SS Рzӆ��	ƚ�{�\B 1�2�X�Xa�`Ӥ��؀��S��7���e� �Q%��X�5�[׈�2bm�ǄQ�f?�����"�M��tğ3��ԁbaG��>�G4[��r����q��7�Ij�t[ۤr�i���H��kC}���K�k������`P�S�0���^��H�q���=�X� �8u�3��S4E� ����_�i'M�6��2���W��xGee�cS��x�FO����@X�v� ��27����$u���Le�����B&>��&���ti�{ho7Q��`�{L�_緤K��|��Zӄ���8�+�]�u��"�=ů�<����N7����x,+'���7��h�f �3�K��;m���ċW�����j��"d���x1�m���$�x̶.e֭'O8��.%(�QW�i���Dl}�d�!d%���3ĒD���=W�.�[v&���Aj����θ�$��͈F (ծcrX,�ĥ�(c�|��#!W�4c�w���&�4|�=@��_�m����x���GcI���"uA�{h�?Q�D� ��,�������B�cPFp�Q+��8�:���r�*�E�[��K#�o����+�<���z���q�muk�Y-�y�����7�
�K��>�2��?���T�jG{i
^v��?�������8��!�{xj������%w�`��WY�8��<�ɜ_gi,����>}*��P����Ya5:����ӳG�t�2�V/��Չ
��u����J����qI�a��?j���f"�ˡ���N;�َ�@'"�_71�;
�z�!eG!ȆA;�O#�����fC�4t���aߐ��;��R<����k�d�-�#S�0���>�6�)��gm�����޷Gݑ�`ڻ�5�����:\��C��&��6Lg��+3�(sc�F���a�$�*{�9���3Gb�<�6�Y�X$ѷ�[�g@�$��>���ß>�[���fVrj���o�#:M�������k�/;��*�KBS���2&�-���#LS�EF	"��4q��Hq�R���� ��s��N�'VG�6=H����H;N��f�!�H��%�W�oH����O�¿Ά�G� �8۾U! VX��.�[>�Ӏ�q������ѫ���N��p�ĜF+@?`�����԰d�L��CԷ�}U P��h�1�[pk�^�,lT�{r�2!�_(��nF�[�x���+B�P������s���(�W%?�����*G'��ޏ�]�
;Z�l&��B�CT�ؑH��09�f��1��ܠu�Ԋ�.���jTϸ�v&��3�/�9>��v�,B���$��d{�Ģ[�dS���<5�#�pf
�x��9���	uO��HH/��H�'���f�E��o��KZb%#�L��9!]r)HP�&2�{� MZ���C3�"2>
݋���y&�˚�'[�f4ݪ�^�ٳ��귻��\��B��R��k"�h�*�/�f�������|��[2pV�5�Z:�����,x��Ƨ��s��Q7 �Uj_M�F̣&vH_C}�'V,1��%�*��enAǛ&��\\�
ՀZ5��<k��l����lB���*�����9�i����{����< P�x�6;F��%�m��e��n/���\u<Lr|�n���_���QY ^����aI��͎�,zz�c&B$6*f�?֪�R�������U��E{,E��';��x���㟋��m>G�	�y*��{ ���S�1��̜�Z����H��3�5��-F���/�E�Em�=p�J2�	A[�2�h�N���_O��#�K1]�I�+Jʍ�E��~ <��r���@A0�p��k<'����~Dl�?HW��?it���_� �F����X&���?�LJb���A7Ϧ�[Z�����h�#Q�̦�l���lU��A�>�����0�?_E'����~��!JDS#�L������u������;�E.����f��#=�%A�o+�G�������;=N`�`�x�#��D��t`(��
��T�@�撺|C=w�q�^�?O�M��nb#��}s`�j��6��:6��"V�u3�2�`(&����쇫ƏR�~�xY�d���C���Ң)��� ����`3��[a��ڦJ�[�@]�و��~��zz��w����ty�nV�����P�v��·h�/ͤ��v����/h |���`#�1������7�dV�+��^���K�����v+���xi����r��P��:04Н�2tF���,���x}��KZ~�$�U�N30[�/<e��_��G�1l�Έ����n�.=��!�������a8����Uf��v~����(L����L�*�ol�1����[��9�+��z����X�H��V]�j��r�Zt�����ҹ���	���9�ﳫ�I�V��,F{1���+_��")�N�i)봅��jqu?�m����g5��~�70(���Sk����O�ޝt��1�Xn��\%������9Gr�Y�i��x}.�!��eW#+k{^�g��F��wu�����v�E����P�w�kv��1�c#�-êL+���I~�=Py������zV���}����*��٪ V��M�=(<�g!�N�s<pb\��X��L��&�['a���i�k̙��RxO�%�������1=����� �l6ϛ0A��wΑ�&G����ۂ�c���vf3�<V����x0�BG�1Z�]X��S(�*� ���Or�6�i:8iz�JJ����.۪n��S��o4]I?L\X����?�<�܅Oc��Q**�R�[cb�?��1��$'�؀Y%��¤o:׻EI�(�M̻�R�X�`��p᭍D\����S�rM���
wwD*���Γt(���>�5�7@q�hO֔��_Po�mxA�|	��#&�*(6�U�[z��:b��ʘrL��;����"��$�p�W��>;<����ps�б�WC�0�0���G�\���=��8ѐ��qd��8�Ǧf3��E[���\���L�+�I3 �^���)��#x\d_���:�N.�?�u��R�c��<�F�X�
kt�~MI���6x/w��Y�uF��`���V���_�k���؄���d�j�xҡ���x�����4�����'֔1!i�x�âiΏ��e'��cl훷H�k
n �>��3��ȑb��
�,p�央WSj:Y1�����kג�uj��4Ξ)!��TzS���˦��*���V��ڌ�����݈ %�D��	�D�Q\�瑕Z�2�v)����#G^�n��� �)��:w|pd*�u�X�#Gv��%�b9NXv{Q�H]��,1���H]ՖR=Vm�{Jd>�k���Gg��>�!-X^Z>aŸ�v�����]É���~uF�ف��D��m�G� 0�|���u�������O(�]��t�r~p�P.�\��O�і҄3<���Bnj4�w~ߟ��,�?[���^�� aW�n�'�獽���B�f���&Р
���y�'��������c��f��N:w�lA̐��P�Ё���ڇ��T��>�	���(y�Q�1�}� SI��{m���=���mٰ2;��FQH�CNK�#�J˄�dÝ����4d�h��]���Hŀ�1̫'n�!M��a�6�1U>W��/��ع�ѕ�?��J�y��hf()���g��ō�0�U�IY�0���B?�ta��:��8C�>��?!zP�u�F��Z�+�&wI��Iu\J���wH=��0W���n��S˶qȪE�`��]9�a`Y���&t�ɿH����d	\x��7�-��u��)��m����A�v������js��Q��X}�g졋A%�Unu+��ҫ8P�v=G�I��q�y�\�J.�|�{2Q3���Y���Nt"1K�b*�1��6nf*_DȆ�d@0�n���ªR�1q� +��$��`���Te
ܕ�ˈ�;!ߝ@�C�җ� �2n���JA�v��u�خ����J^Uڷ�+�����s�X��Z�Ւ5�l��0$_98�I�m�}d�R�]��J��3�!z�g�@�Pg��M����P�m1�.+�'-u�	�����d�H�`A>�#�����7�:�s����vR�"$EG�,�)�"f"��ғ7�I��g:�f�2U��v�����4��g�6%�&ޖ�~U<�?b�r��R�s@t �e� �Y�bS�T.��<�C\�����82��*�c����w��o��	G�����)���w=�7�ļ�K�;LF��rzK��eux�.���|I�i��7��в���t��ʉ*������h1�`�A�,g�+�D�qPx�\��&�1�y�5JSh˃.+JWܙ��ua� ��`��1e���h9&N��M��	�����l�_���?�CTNK�����)n %+u�*o���R�pY��r�W�g��9
����D�%�������T��Q��?����=�'������2�P�\�ׄ�.���H@&Τo7�p3�$���l�,�;-gyubwAHI��ҝ����ݣ����5e� �����)�2㜓�Q�k��
K�/��ܤ�ٯ���clIx=۾W�w`����xR�n�c����\S���9B�/H��ӷtd��?�N�ճ��0��Q���%NT�O�:�R�pM�	j�;t���+����\���&�h�s��R����D����<@4O"��x��ז&j�~џ�mO��z9�j�KdMA@؇������NJdq��z�P�"퀍"���I���c+���*��P?`��]������{�#^�&�Ս\K��l��;���A-�ԝH����Y�\k����_�
�@=ߚN�����.��;���j۞6I��B��R���-�yB�kw9Mj�B��Fʘ�ysm*LB�����z-+l�q��n*�-��J�^���Vٗ�@oƗbb͙�|����H��ig��u׆�����_e��A1�)}�Ĵ�\R��0��:�Ep;�W�yB�{Of�1�t��a1�&Ut�C��la�^�o��r�7^B'��꓾I8qb�����bm�x��E�d��Z�'�+f�}>���ܷ��2b��v��G�V)f�Nd��o*��Wn=�6ZV%�����O2�
W�ߠ��L��IY��jU�N��k]}�׈7iqc�g�.�G����l�Spf��z4�Z~�����]<���ֲ0��^�A�Ӏo�㕯Ğn��nme��@x�g��2 ��_%��\�J{�ڵ�8u�4�W~��5<�:�d��9~"��;��m=����!/�qVN��I�e���THG!�����}۔���2N?
�����@�J������U����w8�̖�gKb_e��:�������q;8Bp��37D�!���OyII���c��E�qjnm>�:J>8Ӟ[�Y�����0��n��f���4z� 4.�$)a�J��)���胣�F��Q�	_�����k_������{T�x�y�������jK>U��;��e{ 5­��S~4R���Õ�%���N��Q�[�7���R)GG�������ր��o�Q�!��y:�=�ԡ��n6^ZH��>��V#
ݑ��c�}+��I�ݎ���[��"��4�_�^`��Þ�}����^B�����P�gL�������gf=(�BU�tkK	��O�������1[!�K��m������������|*�;M�ɘ��D�-R$���-�s]&V$�>�+���������&�C�(�N}��^�I.qD�kj&$c�#o3�T-���;��h1�������)��!W�la��i8f��.S	�vNd�,K�����ю������|Ej���$滺�����i6��a�JX�K�J8��H�kM~�P�����Gȑ?�'���˲MA;��'�]%�Hkh�=�ɨ\^�s4��� 4_�"��̈́��Y$�٣y=�����~W�d�t��
�8�2���rh$�٘.�O�N���%7Ψ�[*�J��h�y�Q
�e$���I�*o�^h�u9M��H�ΛKx���^��mw��?KT�'��p�t���	^xW!��QC�v,��%{�[�ťc��x��?����
d΢u阞��l��wb����N7+!�
��'�T�%(�/���b����/�Xg�a�U!4�-��
t�0�{3v�֦4��h��VW��N^��2O�%y�ɂ$���3�y���7ӯ��ay�M��aM��2��~�(C�ȆË�݁7M�7l�O��xMƓsǗO�^ΰ����2I�)���ڡ�XV��t�p�
�2����KC)NIOŅ/�y()��G���wJ�/� ����ʿl)b�#C�Mݻ�ce-��/��@7�[x�-����T�'=�RF1s��ͯp������h-�E��Z�����nMg�-����S6�ώj�#$���K�g�N�f:�J���΅���E/���y����j�~_0O���v��.B1��~�]��B�u� :�(�Q�� ��?�"�׹�E�z�*���f�Z�LD�����ne�q4��e_�@���w��� .yzI��h�_���]�B^�<�#,��1W̹��'ے�N��qI��*��D�����h�s��	�����G6!1��)����!Ro�! Ǽs��Ym	�P?z_�P�V���%���u����`�-��)B�8!Hkc��9�| �F�Gx�:��t9fF��Oi�xs�L[]3��Z9��ՑNq
�`q�I�r�e�������lX{}�3}o0d-�D�Lb�W�G�x VB�H�xH�������&$f�i}I�[R�bxƜ��S�{B�>p.�){����Kq�?���] I�޸��v�Х����G���l
N�n�@w���HR��Ν�'=tu�)��lF>��oLu[W��M���%6��E-�B�	v��G��}���җ?�H֩������[��y;�D�aYY���:����T�L�B��-�#m�sڸ&��V�v���R�,7��������k#V��!�eTuQ��T�	v n3;i�]�©%FV�� �&/_<���:No`:GI����3�Sj��P7z���#Q�왨��;�Wf��Z����$�f��%�c��6�5 ����y�ȹ�H�r��1玠���HYG
KP�(m�nP�ck̮�H��%��PI��G�g�����3k����{z�0�����t�Id�K$]��W������Ne�.X=hI�����0��O%%`�qV�TR������/-}��<z���ï�^85��6A���g1�Q��P;��_�'8B|#�-�iWRbKkh��=�`T��H
&�?�&�0�{�%g�"~��Ƨ�d0����f�f��B���NO��蛋��$Q�l�d��LN�v�sCB���2W�J�;v���.���!��/��&��,ӣ~�	��4�4�)��f��3FR�蚻GT�5��z����1z�Fjk�f��vw&��F�OV-��^:�
{�u2�l@�����{�7��[��*4�e���A��ԇ�5Q��%n2����P�����s끏��
S��R�X�{�e!N�{x���>���d�S9*�PB�I�EL�b�r���C��g�M����K�G����a6�.��"~%�O��'��+$OI�_��#��A�H=�t����|3c�лzB*�i�A������A�g�|���1nUٶM���d��F/=�Wc+�I��̌h�\Ҁ~ %~�)�B3�%�/��pp[e�	QC`��(�(��a�L'�wU�M4\�d \������v��-C���^�v.}q�ǧre sG;\��:E�yᤔ����X�3EpM3�h` ]&�!���^61$'�P�@`GvɠϺ1��m0p�����"��V�,:F?�f�t�'^L�"*q�o����Kz���=�}��lJ�dIr�����qj�w¨�w�"�<VS��ٌ�M�q�K�:q%�_ �ܵ��.&)���P��,�(�[�l����U�a���8�D�U	���R��4L�
�ӈ��3�/t�0M*Ѫvl�RUN,�u_$����_��{r�G�T%ZW�U3��"wߚ$ !�V���ʋ���Җ5i��涾�w)���S�
T)#�%�=B�р�z0�ceв7,��\�C���lM���6�_�eM1^�#Y��1�?HAG��b5:�563@�,ݎ�`2a����?�,$7&�8a�z�R,�%�>�:�PZ
���8w!bm�l�4	���}y�#?�%B6�c�^��7��!_m9����DGP��-��"�ԍ1e����!#5 �\&����;t9{��K;��Y3B?8�D�V��.v�'���ي٤���=��2-���;џ�L/�_�9|����P�;=��7��L��s�}���V�U.."9��7��2�5w=�˕�������-fe"�������{���e�-]�"�IW��%�}8(Q�8������_����R)}�|z|&<���6%���
���6��:����d᭘ j�
U�|,�n�9�Š��oE���|�]�9EVg�*IF9���'e?^;�_��	� ���I��}��:�ѿO�u"�DA2��a��x��Q�XΏ��@���s"� e<4N���'���TXB�z!d���ʋ�?���(+�plg[ۺC1v���-Ӆ�=	P�c�!�_�)���
4�aZ�/^ަ���IT�����;,�q���2���$��x�!9n����Y"�6�[BDoWf]&�|
J���}��/������Z<K��Q5W��Jǈ:�hr��.���w��7�t$�d+�KR�Ά.��L�n�y����/��M�^x�B����E�_[5��M��I��vf2]=�Jv}��!��!}��X�=˲�~�eJi��Х �U˓�aeU̚����
����h<��K��.9:����3�9<>�3[x^~-}�od���	oř�!z&�������5�Rw1����浐�,�ʖPF�o��?��	�[$��2�K�C�D����i�[��b��|݌��r�^��G� ޵�t_��Ij���k)t�/�$(�A�����X�U�<�����4q��9���Wh�r����\���vS�os�n�T@��/;�9r�J���kpb�<�dД��F7��sȍH]Y�"בT�1��\?��V�K�0d�`݋�%i�[̍�)��}+��i!D�`꒢~z��� ��ڭߏdq/Y���6Sa=�h��H��=��� -���l��(v:��Q���+a�4���i[����`���x�Q�?,{šo#�/ f��]���h+����N	O�hne,�R������m��yZ={�.wrDZ���>.�'8��+���� ^2��/	�0���fz��L��a��{o��vڎ'e� ��� ����::�J�qAb�����Ү�$�_�g��iW�n��B��;6�i��|)6�6��"��E�=����d�]���4�.H� f�0Ti�V�"�gnM:XFw	fןe� W�%	{x�t5�]�ٓc��Ʉ�=\�ӹ��5�����"��L�a����J��W���"�@���g�'>&�6��w���8�:��������\�7-����[�Pd8���Q̧��%�u��^{�c������a j�xoU�a9Y+QT���uCG�f������Q$;��}��BQޛg�։j�^>��C(4j[q-�����;u�`�=m�	t+j�:��3^YP�}2ƏHH��������1����}U�.O�A�=u)t'�$P!T�Be�5����`�5;��j�ﭠ��
��_��U~�.r �(3L柢XRY�
҇P���\0	c !�+]��JQ��6��>q-�:�7�2/S��L�Qe}�P��rN���^���ީ.�54<F��� @s`�R�����,�\p�A��
��[Ԕ���Ƿ[�A�����!ͯ�ݼ)0���D��t����y��z�@(s!  3W���C��r*w��T�Mc��� D] �IUr�Z3Te!Rv�ɏ�=V^����	����C���(�?��� �lk�B?\ma��^��� �~��&��[���>���!���ׅ~���J��7n�
�ف����Q_0Zcr�[�� �1�%��9]3V�t�/{�U���?GUJ��ئT�4��}F_om9���l���>X�t����1FwY��t�<��4�Pa�� �uU\��(JQ,��j��E��,@޵aW���O�Nn�^�9#� LrkfC��++�g�#���T��z��%�-K�4�6�����|�����HI�Y����O}���K��I6Cˁ6%bK~�1�H+M����, j�1�K\��n?Bw�O&foT���x��B���Ҭ�؟�,���/,w>�a�3^���L��N,D�ۖU�e�;���Ƣ��	�QI�2�����w���EL����R�C�5�[�io&Y1�M����9�k74�*֫�b7'����ᱨD������A��=��!0����ps���YGSa�Z���>R�L��v6B����4<���zm�e`�%��e����['��(�d��Y8tsų��7h��ك�󆠷ffA[t}�X&�B
��G
��k�������GfB����B�^�[F�\��U���yg�C��ݯg�h!j�� Ծ$�
hyP���ZN8��Jz��.(hй������2��3GC.�>������B1��N BR�O8�P�h�L�n�R̘@���:���F���96��HP:zwQ���V���:��+{������dzSw������@���U�]7�[ax����sI�� �X�|�۪Qyݻ_�@�z�ȓ����D7D8F��a��ڹ350��7&@<�5�g��{�H
8'v�د-.�mj_g��]Sѹ��҂V�y:(;�O۶<�ѯ/䬘n��xd��I?�m7_�Y9[[�	B6�;4R�|��n����-��~[�����=�K���t;� �'[S�#��M,���Ue΋ʷ��6����go��<ٟE�觶B7UBɎA��߷>>w	by����	�i�����J�����ܖKwE�y$jxs��U'��jJ�0�Ye�yƝM ��=tg}�lJ���GL��:���N2ؽ�roՏ�XA��W�U�~��	�M�K.���{:[	�u˿�@���k�Rzx�2T���hJӉ�U��r2@),��$0Ç�k���=h�߹�G���ø$�ʇ�ФB���>�O�V�����L���Q���8rG2�>H�H6�����8�f�fu��lN��*�get��f��y�uﱣ]g�m�9fn���l�Hz�D�b4';�\���Ԫ�@���g3E�M�GFC2B4�4Iy�;���+3�BK-^��*T�7��GKN^�8\��ib��t��@Z�#eJ�t��ǐ�;,�gO3}�g�݇��~�1�|_��v(�sU;�|��Y1��C�U�}k*�x�����ƝeH$+����k��Ӷ�5��%�.+}ɬ�z�F���1Fm}i�!�w�'�}�q��.|���GI�n'B����$���5!�=�w���G[��EF�@��S�[R�O����r�����q�M͂&t��kd�L�����TW��BFJqx�l*��  ILCP)=���qYLYJ����hY�Bp�bP4���<���C)W�� ��edv�p�K�kU���n\����.d����V�Ik�R��4�:hb>��Eǫ7�����ջCe�N�bO�H�˴h��2��U;O��*�|z����w]f��KMH,-��ڑ�q;,�=�Ed�E�o׉��O{���#��b��PC��,��ĕ�&]�GϪ�"g�S Q'�نm�Й�GD�X��O�#C��m������Z��p���J�UM�j�����7"�7y{�R�����P�����0�Y3/L�솒�[��X~�M�\0t�t����@�c� �U��.�&�ۣ*����Py���R�ez}���1m\��*���B؀���5�U���(�H����0�xW(⢃[.<�*�D"q�cU��.�����D����L45���� C���a���355unx7��ބ�9����	8_�C(×��>�8uW^�*�@��{�GR�$²7X��׵��!���2���;n���+��L��<I�!(�{�����y���<9Wz�[�Vh�@C��Ya�����"dn���~6w'�D�A�㇬v?ޠ'��dB�Bu�w�kP�G���fN��(EdK����(ģڠ:��/�E�=����/�Ӷw�@���eb<,hQ�*�{`�=Qm�b������vE�-^w҃�*���T?I4�в����q�����M�	:��6�������ĺk����W�1���\/"rփ�YU�Հ�(]�NS�e�����U~�PI/��.��N��$ί��(��(,#�Ѝ@�O (r��5�7�0���Ƿ�t�p9ݏ�k��
˕�[�{�Z���J5O�嬒�)W����ɈM<x
���o��iЮԓ̯�����B��� �p	0�F)E����*����1|�@���E�}7�?���+�M����
���-�,���G�!зa�U+�myvg�B�q��k\�! C��)@�0|�-_���V:���m��(�ϱ��h�߆�ֱaQ(�2���4�7�lzH��X�v���rR��w�B��2�JOѻ �*�"��Aa-ɢ'Mxu���Mi-]uߦ�����e�]����^�qW����Lj�@��4�.�5�+c�X�tV����X�:R�Y�z���<b�����R�N�0�e���?�]�ʷ�摬�3=��J����������Y�Oܼ!'tg#â���:
�qQHdC��;�f�Y�I��c���꺈��l�V��Ӷ���'Q,�d!vz��:C�����2�.��`��#����У��z�l�Z�Á�$��x���+E����Ǐ�5v�L(8Du�s�p7]�&h��$8����(�"�V�Tᔣ7�F��/0����ֱًS�!q-��v�>7��.��� �5�iIg�Ӭ������Z8ˋܵ��rQ��7�fGg�:�<mK�D�M�V)c
y�Z)��D��iq�`�Ma�)�h^´ge��W��R*���J�y_i��ؚ�dT�DCS����?i"�[a~���ΰ�S2��Jd��	4^�A��߸�؃v��D3�7'n3 5��Q�r�d�ߞ��lr�4�=F+�+�������8�F!�],��O��nd�B��A�����k��w�Ю4�$x:U�d��Dh$��jm�OD���.�:`^�8+ϲ���<Y�ٵP/�X����¤�v��ށ��t�E#Ti�6Q�����2����7ͳ��-_���|K+�� ,Ѻ���F|�1��Kd�61k��{"'#x��T3AQ�ղ}J2R���=N��c�LZ�Nh����r��S�_b�'�(T�K�����8׾[�@�f`0ʹ��|�(��)l뉱i�Jl�����H/��'P���Ju�����b�nQt����O(����p��y1p����*~CmEiX����qzK��6��v*��h���9D{��Ȳ�EY�oVYj��oM�Bq�<�C�Ɗ��f�6xGrw}�S��l�@�6<fCU̿tζ��CW���`"6�ƽŐ&ew�V�E?�Z�r`�y���Ud~M��L3��k%f��Zظ�R��T"�`��$��͑��1��6�:��t4��%��J�x���pW�dv�qlԷ���OٲF�k����+�?�(��t�������QU!z���r?:-t|�މ��h`�d�	@��Abm�s�%�d�U��X��u�C�w�[t2S���P7�@^���+��7��!�w_0�w����������-�s)���=�7�2/����%�m����d�QɊ�_ʻ���I�`�"�(`�S���u���9�.��
9u7��.dr�Q0�P�$27	���P8a~����Y�s˂?����t��X�n�ڹ�u |_���>&�7��
V���w�8� �fCpqD�J���!�zAE�n9hjDTWѣ�+�E�j��s���g�T~ ����%@2�t��(����D�<W������]�]�~lv��b`���ܘ-�&��}z���vȟ��0�����.�֝a����Ώ�ʻ�G�,Ks��HN�3��3D���E8�����~�)�)R3�R� 	8��0��7;r��Uݲv;O���(i� De��74m9YQr�J��01��57��ު^ ����ߪ�~��B�ɮ�9�\M@U��#S ����H�t��@�U�/�yI���䁞vR�y�z��~�YB�
�����xCp�ǾB�M�M��UBk����z0v���?�w������m;��볘9�V�E�N2��wvA�R����a��f^ظ����H��˂�1m�9ҀK��{�W��j��9R�'	s`�F��L��K5ݲ�W�h������?K織�Ô���tK�տ$w1���2�)� �6�$řW8g��J@�Z|��0g;]M�h�g6�\eemNs���.[����h�?����t+wM��� �ey�����&����b�_[Á��	�?{k3�T�tU�ty)�v��;���e! �DD3ulny�f��݁L_�H�=�/�o�ŗf�rěc,`v`��7	}��蚴o�ۖ/$�A墨�i�WZ���f|�j?�����Mn�S,x7O�^��~Y߳��RFok��ӝݽ�(B�\H�{m��M�.Z`� Nv�K9�L�T,b��Ex�o�t�ۓƴl�&�峉<a�?�O��'�^a}oֳN��qm\֚�f%!���>��y��k�1�yn5�J�0$�l�A��c�o]t��Q#�I�7�;f�&�����B����3k)�ZįK�z<��lV�������9�ߛG>������ԣ�oȟ8��؛?ԍ,�\����.�ӑ��X�@L]a`-|�E�� ���Ǒ2wb�"����Ί$[֓���P *\�+*"�Y�}��#�.�g��-�8\��t��1K�[�)�Hߘh�� �ip����Ch�A�\�d9��+�z�7�~��o�,��5��*Ŧ���v�d��&@��pd��eI����pw=�^D�-:�@�=�#���Բ��
6J��X�#_,�(~r@\�NXxh�ѥ8��;�w⏡ڒ	b�D�R�Yz,�ˬ.���`�.�r�bο(��K$���"�y�#� ��VJ��`ƈ�{�ؓ��Y0�y֤�W���W��]�)��[��u��.ş��<ˈM�l��Qg��T/���͚�  9
3,E�٤q�a���ouy�[�l?��}������P܁ګ�tx���V���!�˸q0����!��㮃���ߊ{+h|�5�n�L�r�����F ���������~Yu҈�o!�����2��0��*�Rg`'zsk����e[�`E���U��h��[�)�o�b!'���S��?tQ{��� PǜtQȱQȣ�e}�$�eHT�(���P۲T�����`:�W��ު�7[+�Y�	u	�U@�N��ˊ�a�w�)���k�d�]9��N+�c��Fj/��{(��	����ODf>Ō �����Z+up�%��{�u�ec�Ui�%j۴�|s:e�r~�hIF~����y�Ӆ�Y��0(��Yi��;Kr�(ɛ�(_隝C,�k$�	f>�P�X�����`�}m}-12hIB��Es� Q��.�%���Wi;��Q�a3~S�]Ǆj@��n�Ԕ7��|�GzeRa~lxb�W��ǦTV":�l
���A�=~���(�(dD��䉚�^�u_I0�m�����6N\&��(��@�u`�`E�����g�:,�F�H�9����u�j�.v|�;@+��&�I�\396�Wv2���IS'��d���9E�yf�]�$���.8�f�Ɠ�?uO`��@o�D�ga���k��b�ߗ�e�?����v%r}�Q���|�ja�.�e� �M��>��yI�����p�v�M,���L�I��B*�x�L�D�kh�Ӿ7���ƏoЩ^�S>rqb3���<e}�o��4�ڻY�N�Ϩ*Q�w�eZii��x����Qaf�5R�1��n�J���l��G�}o���I�8����dE-�Z�2��X��V����B54����@��#�6�*o��d'�޼���{�)k'(��j��^s��)�$�,.�^ X�p?N��k�!��g�T��)�~1uU�a�}�AxO��"㛊���3Y��<Ȯg�!�k����8i��9����]d�V�]<�3���^�-1������tל���y.�dA���"���Ш�%�2���Y�9N
���`�;�2��7;���[�I7rU��P�������U)	�� E1���z=���rTj��;�)ƃ�h����uj&��@�Hȫ
�B0p��3���Ɩ��Z�) �ϫ�^��lw�זû'�*q����`�c��/��
�[)�7�5��L<~��D0�����0(!ӞB��-l�F����յ@�P�ICǟ3Fa��o[�Bi�����Q���21�@GKz�b�p?sԅU#��:��V���E�N��s��ks}��7ȺL/��ƌ��(��Κ�/֮�ǡB	��R<�}��!OCEp�Xa����b�0[TŘICB1:w��r]S�C�Z��~�b��ǋׂv������ܿ�by���pkp0Er�=��w��O(ay��dX��fo!J��;�i��#Z�1��H���ڀ�$*B�vR(�Q�����M�W�:1��w��]dޱ7ЕԿ�-���k�v�k,6�]��sJԯ���r���	A����e�3�}�A#;�!̝XUlh���)aCڃ��i�4l��i�UQ���/W�	��A�A#�!�Ӱ���6?×xTx�	Z���MG�8-��K���ٹ� ��,5�f�2�D_���y+� S��ʩG��g�/,̝��4\M�t���&AYM蒲��]Ʌ�<�Ĝ9:��my�kC��G�.ۏ��������3�R�q�٢���?�Z�wE=`��S�0h������3��F�z�M:���w�;`%2bM��M�D������v���/��V$NL�E5�$A_ؼ�/J����^#N"���td������ei_���,��d���e������N$������G#� �o��	H9��"�C�̠�]�K�2��4K���r9%�
O
��*����za�Z!j�=C�q=f{kڀ��jMb���wʨ��fB
�5���l�ϔL_��;���{XL\ͩf�����çzR�&~�5�=M�/I�͛�XA�O��&Y4�����KG�9d�$��P�-j}�K�g�*mX mAį�� ������"����#�%}��+��a��T6m1���;^�h#�g�V!���R>��;�xk��c�A��H�U��eK0	���ox�;Ķ�ހ?����&��*OVk�RUv|������e�HS΄�&Tr���m�ƱUW�i�pРRwv��<�w�i����|�W�$3�:e@D�
>-��r�u�������3x�!g5[k��UkD�@�3���<�����A�F{y���FH�t�W��/�S�Bߌ��>�wA�p�Z�ѥ���_>O\[oq�5S�5sX��@i�m�W�m[�o#n.�н�Ʀ�H���^ZC������߯ ��"��+����7H[
�.�+}7B�<�P"&C�#�{��RL�d�E{؆�Q��f�Ey`9�l��g;U��!���lw6)k���V?y|��@�6(�/y���3��;�G�/W�J�@���O�]	K�3���Q�����꣒�o��߇*QO���)���vCU�E�Ï��IZ��s�$�b��d�o��#=͓�·���,�e�?h3N�,�#O���!y�xmc/�x⟌^`2ڴ����'���q5+xE�Wtֺ׸���H��� �%��0}H?��g*�kN� �������f����^.����b�ۂ�g�l#^���H%�ܘ�*u�&��j>�3���0|^|�QP"��
<��i;7���K۱�9[S�ɚ�̖��!P�X���ڴ�� zO�]����������8�=*��Lu�0�5-
��6lL��)�.�&K������?�x�f��A�ʉ��lE�I��ɫ��|�c�p��
��9�H�.�⥓hA��ic���Pa����tm�4��4Ɑh0z3>���覞���d��0H��|��,�Wj
�W%d8�F�c�'���iI�<.RZ&6bYx��w���G���q��fO�5�`�D(�C�l�T�ZͰY)�D��%�{T�_C�7`!�Ƴ�������$彨���oVVΆW�? /٨+��tf��eA�
�����c�-��Xz�ڀ����׹�#�P�W��3,���Tt���ۥ�d�����P��o�A+���VO�G.�T���҉#��G\^����3T�!W7S�9�U+�����.�,7�Sa��[��r��� f�"6UV%�&���Q���Ǚ�:ꏶ*�Z\�\b�Ň�9��A���87QzwC�ʆk���>��Ug�3/�D#@�w��[ԡ�	Y"���_t��ֽ���+	�O�� A����n�s8c�v�rgv���q<���$���/?��R��
��ސ���R�X�A���c����+� ���&�S��[M��yrji�d�	p�@y�s�5^�p�Z� B�!1��Ak8����?<�qZ���}���v~��-_��#�5��s��V~���Ī�5(����5��������kJ�,F�NW5f�D9���o�f5)��93��0]c=�G��Y�O�<[9s^�l47�$D�*n/�[��M-@g�c�BސDT��xE
����!�/�����b�_������`=2Q�������D5*�(P��B"4.�c8���%��@�+���tȓ��${p���6;h �V۱�%�g�["�^
�_���,j_Y�ЅNg�(6E.��P��s1!TSh^W���F[�,���f���Ui� N�2ݳ7�o��ŗ��y�m^#�Q�1���u��h�4I�0���H�Ī#K|��"z���8��UY��YF�F�^lV|���=ϰ?�Q��� Id"�b�(A���H)8��aCG��wS�_�!e(+�2�r�`��v����F����������z�.�;����+���9��@�ZK6���C�����l}�L�����c=_P_��*����ܤN֗�"A�}Q3�F���XlzUAv��X#��z+$�M0<��+9�[�����<l�${C����͌�'����璕�(c���"Eb�д�r��}���y0�� vj���G��>
=Kw�: �bd��n[\+���W�j�+��uSAG]l�W��鉣�ݥ�h=��
�n�e�����_CY���&�I���̯�`����)}+�J���:m)�d�~8S�����v��`o���ʺ�'Ψ�0\ uTI�i�yy�P��!�˵HA�@c�-��H��*�*=��0�A��`l��6�A��R�k�Zdeps�E�Ա~��r�c�ຟ.D�VB��'2�NO^���G
��?
��7a-�_�+W�;��	���T�)��YD���R���ڇ��Ҭ� �3H@B�-�-��L���MpHf-K}���}�c�ؚ �0+H��A�l���Τ��r�@��A��Z�GjգR�5/ �/_I�ZS�2�|`��Q%�]�2��h9l�ȲIdeT��������/jY�K��3��Ƽ���R��J��(8�Ыˣ�$�Eo�n
^�i=������_
��n���8�h6�V��O����};Ը[5���n�%�eq�V��$M�ڽD����:���}��I��Ϯ�f[V��F�_$�	:��c�.�7���nk	��	Cn�HQ���~f;�^�����Zҧ�(�c�`��;�C�)���p��&��O����ܡ䖸����
�#�F����sN�g/{��L&�Fe��^2��� �_vuw	#�lC
�bKb�gJ�+b���QL�[��f�l�U�>���r�͖�*x�Mז¯�$dep��Z�z��b�^>�"~u9��u�;bo-{����Fw��U��ę�G��b�Й��60�u���#1Tz<��A����H�V1L$�),7��K6�e-]A����{��-ت�����T��^0�m�%fD�7�}"XdZ^������r�����A���C�:PNh�'�hq[c(#~�f[peI>a\���FYG�{��W�)��oă�R
�S��{1�����M4�z��`RWE�E�m^�AR�į��|�k�._3tB�A�6i�����&�|=o���0^ӟ���i���`���}m���&F��-�\�A�j~�M����A�a��K����1S�Ӝ8�XJb�ϱ����=�ϡ%_p�.���I����8����[��>{�o�d{�^]���;Z�x3��0���>��!Gzj	��EjJz3�ЭB�73+{�F���R{�s���_
�gV�F%��s��ů �p����*�����q}��j�n�/
+D3�b�Y�o�����t9�@'�<�[b@���*����O�3��<���?�f�e�vZ�,6�HH|P-�!!�!�����|��:�y�Ї��� NGV9��cV���vG��v&w�Iv���F�.�]�X]O��팠:�����
�ӳ��{o��6�_�5��]�����!h5.�O�S�����U "����D�}-�{¦�C��$)�#��*n�,�O4�~K��G<�X,���OC"��S'fm� ����8�]�E����_jb��C������"c>qo/m{�I�>�B��m\�۫b`����� UO�����ն��S6J�JP`M������V���%z��l�+�U������O���Nf�w�������zP'�6��� ��N�s�����U0\�b��Ee٣N}�c/�]|&�a�B�*�UM�t��lG������p������l�����o���%+}B��d�BrG���Hi�X�bA���7���t_�m���J+����x��tY����M�kq%J���5����s�w���� �w�rQ����FO��_�|��y�qڨ�&k�׾�B�c�����x��"�ٵ^1��4�٬�A�"�O�b���,��������-W����V�M���1Л�8��r���5Mb߾a�"Q�)�Q��|D���U��q�k%�|��~����W���%���A����
#0!Ͷ>.��YE�_+�'ccpaPO�Α�x���.=C|I�$�������a��������2M��f �!p�`��%w R��t!���@P�s7�
-o]f_J�&O��R{�ky/u$/��} �F�qS����;d���$p
d0��D��Yj�\�'p��7�ZŰ)��%Q$���(X��-?���nWgxN����}��{#�	�M1z�������y�+8��t ���Q*��1�v����d�!���h�]V�q�����=�5�m $�'S���ⶻ�'vMB}�rw} ��A����R�QN�]d�����<��7�(�#��σ��o�+�U�^3�澵�
��֫ ���2{�ܫ��YC'�F۞�v�`�|��b�. ���1&�����x���Wl�	��C*;J��cU�nM@�s�iG���e+��i�H���SV�3�@�.	c,7�[��]�k��VV�]U3�ý�fR����؅�_t͆Dg�^2Iq�����f�=�X�ij`A`͉�H�3�I��E«nܵE{�݂gO0}ג���꘹�<�C����p&���ߺ�,�s�n�t�3)	��g,+�Sa�+)w��$��Se��F�
B�+�b^�]�g/V�e�m(��-�xGVL���*���b�Q|9��?�3#;�Rd����_܋����Hֻ�
�n�z��<�u��Q���`�K�3gz�� u��>�L�{2`8v����i*��0P�i{�Ԡ^���K�X����!����g��'�jy�D��ޭ��"Z������-˔w�Y ��� pÓ\ں��&���Y{�]�	=�J��oG|��;t��<\�ԧC���Z��M?°�@���>6�^3P9$	t:�'�:��WMmP}*��md9d(��:�R&?W�XD��OzTY��r�I7��1fV���?a�;���04:��mY��pf/�:K;�?���v��� �?�	�i�i����5]oK ���J�Q���vD�*��
\�*VM����}u�л�,;�x��C�I�)��0��m5U�̑�������T&k��P��;Ϝ��0�C�$�#H�&ed�Rm��{8�����O�)�5����9F��d��@q��7%��,]w��z_�=���]�%e���ATmNᛁ�����̻Zg^m����D����j9q589�Y1���'�y�5������H��Q�H�HG[ �ӌ�.��	���Ho�vR���6j���uxh
�0˳z�ݕ�o�/T��'2�r�� F�7�8f�����Mpޤ�!%�t�HNF@?7�KZ��q8�H�o��|�+�Q��Xy��F����K
�N�R�+����K�b�¦C�n���,�K]��T�A��Y��^��ʸ���[�e��a�8�႞\��jE�,~�P7�&�r2���%�r�"q�����!�cbw:#�㺌��&$���>�L�9�����Srե���"@���
��=�D�����5s�eZ���uk�L��蒜��lG{��5�M�)���$m����9M�U��"��a��_�
E|F�z-���Gw��'�Ͳ�i;�j^�D(G�,�<�C����w�U%o	���G={�� ��q��T�7jtW�pdh9�'|ۉ99�[�2/�͟�UT�	�xhT��J��?Oz�Pu)O��$m� ���7������������66�4��/[�A��`�ҙѥ��K�Z�����&u�H���癀�u!�Fk%��/�T&��T.�:��W��ʌ)�`���h���w4ʺ! �xWϳ]"�F!7�?��·i=3�d�;:p
{�B�_�K��
dd��my���QzsS4 y�����;Li�ɛ��Ȯ��h�c���H�.��"�6W�4v�	9x��9����i������^:��LA��H����F��n��ޫCřR�,������|��E��*��H��i��~�o�KA�&m����?�o������Bx �O�3�"%�Hm���{�oW�Ѷ\W�	H/|g���)�tMalM�f��e�=Q$�~B�ds����%:9��� E�R�S}�B~�<�ڳ�C�v8ٲ.���|�g��m�F�<��1q|�d���,� j�E�	9A�R����/j��]�`g��5�V�;���V�[Ee�*�=ee�ҳ��&|i\�qo� ����sB���5|�Ã��x�P�q��)009��R�
��cpJ��QF��E���FθG�7p�t��K�F!x
8MU
�&Y�����#~Wt����ޞW���{k}��,�9��i������'��UKl�"�0����3�3�*̼�ɡ�J�v�N�j/�"��7i��o
G�@u�5X�Z�kf��5}��!BH���������
���T�s����$kیJ��~b�;`X??1,��pd�w��Rw~�T��y���/�ŞI�j��y�=g�zizd����O��gT�W2	�N�4�2w,[r�;�Ga{����diy}º��<�#�5���sX+b�����M\G�^�-�!8 �{�kX�m	�1��иތ�L��.�Wx�#zBMCK�A�-���Vq�`�G���x�����#G_����h��:��~���_=���T@0�-��a��՛�D�5���`jr�RYVt;���e0Z��Q�ګ���>�k���Op�\g�9\Vz��&)6�����:�m�N�x^	I���v���Nc�a��ʌo�Q��l70II�w����o��*���5�ߪt[pw����zH�^5WF߭ R��b�J�[`9t9��b ̑��ڣ}��U�tz��Ƨ/�Gׂ��n1 �O��y��SSE��zA��`7f�@�'4#HY���AQ���� ��{�
:� )77��E-�ke ቪ{*ƿ���?l��@����gle��� ��v�^��*Ac ��*'����yjv?�͡8�׮�k	�"���[�)3Y����)���C���w�,�8�(X�քj ��� Ow�匘�<Y)���aNS�n���`7�ws�i�P��}��c��T_|h������`�=s��ZW�&ΧV�{3p�}�(K�'������������{�W�X�nTLLw���I�
�w��E���Ɉہ�$9|�d�̱Qs�pB��MUN�O{�e�"�?�̭�n��V̱��<e�d�nϰ������w1et'�""�H(��*����L7O�-Z�����a�Y�� �'X�^��{(;��&TLc��[�A������ 5�a������Ui���[[�&���dQ{����c�L^j	�Z��F.�g��<_��yh���%�!������f�yB��:�~��:I7��+Ŷ���	��˷���E�a�H���-���ԟ,�%u��F���j�rm��
F$e�+�� i��L��'��#�O�	2��to覄��T�����H���uԨ`T����z 0��PEI���	fZW�6�S���7Vk�i�E�Ka1�t��!mK7:�chۿ-��5Wx'��v���&��q+t�g�H���������5��ut�׹�h�+���,����GL�G
sَ�ns���*蓚�\-�\�er����y�����`�ڠ���I7��v���^y�����6E�Z�-������ؕsa���Gg�˸�<Ҥ�����[3����Ow��Ldڂ�/F��^�ޒa�#aĜ"Y��ɥ	�1g醍�-��\9ؑ%j�Ɖ��o�I	у�$��$�p S�Lea ����<3���_ ��lz��L*"�׽]���f|2�;^��Ԇ5��#n��b�0�f��'bVV$����<~�;ʹ�e�=VP�Op=#k�A�
���!&���)2�D���8Z�c�t�ٰ[��V
G�a�[�C@�uV�&�~u�Z|kHå�=����Ezݥ9(�e�%Ds�;E���*:��^Mֿo9(���l������N�IM�l����C���ض�$���kS�VV��qz���4jh���>��%���O�����Ŀph���fM����ݑ~�D����.���;�{y��)_�����T�~
b�w5;����Z����В�JVs����lhgj��H�-��;��8�U^v�Q_�߅fs��N����<�L�:dKrB����&Y��;{������>n��ן��¦'}�&y��-^y0q&�٩MC�m�h�8u��)	��FACPB�BT�C^���J�ep�c����h��/-M���9�a�����(�F����/�3_kg�m�0� �Aݩ����m��&��]�AN!%l�`���%�/ۓb	��+�����oL�}o�'kt�s�B�<�?&nhN }��Na�3����,HE��5O�nI�5F�����d��k�$m���Pk%!�W&�����V�a�^"���~���<���v�$�c +5l��^��&Tk�ԙz��Y��j��
Ǘ3��=� �f�.�yw��>�;�����cM���ZȲU�NQ�.�a��A'I���'׏��ˡ��	��1�E�}߆������>��ϟ'�"���>Gʉ���]�-�Ǹ4)��I8R�xgh��o	�Ӏ��u�է��N��1�/X8@|E��e�1�f�H"��1���_�??rS2C�/��f𐜍~u��(G�A넻x�����q�J������6&�$�A�m�N ����j�G;�R4��X��t%z�.z�����z��F�{��C��݂���Λt|/(5���m�*�0.��V�[�� G�4�R~>��u��ۦ��z�r0X¶�"�eG���ӈ?���':5h8�k� �V��]���l�>t&w�6fY8[�#�ia~Թ-�壹0pXs.!)Of��+���eʭ�4����P��r<�z�Gw�O�V++:V�0�\a��E�UC	��;�t�Ǟ�J$V����Δ�(W�%Q�ٗh�\ZB^�b���E%�
�r�D��f�0"|Y��3�~��F�o�ź(�}P.!��q��hp��r�t�_?��Wʞ��شn�{�g�������h��&�Ϭ��y�id�cVS�/krWg&S��nv┞�~��_`�eu��gI���j`� R�ެ�ur���E9E?���|\Л$�E�X�Ê�aaYm��� QF���"|s���I���,�w���g�樔���䘦�U%߱DjO� ����.�{~A���>(�X���m5�\�lp�� !�5��0�"�u�΁x�~tv����-/����3pA�U�iMU]�:�X���w�+���Ix�6v$�q�W�-o��;DB�Z�P�$-��^�H�y��9�8�\&���&��� �΀�jY��(#���
���}��}��	 9�d6�T�:�� ��^�ҞV"	m'F	�c�F�$.�*�v�Ͳ1�&<��/K�7�!�v�&������t �D
�Y�6wU����LH��c���O��Q�37zꈞ'�r	 �Y35��xRv������8��<o�DAM8c�1�e�@@1���)�"�;p3�e6&���:�(�5^��9n1Xbҙ���u��XCG*J �i�A�k�P��أ�\<�?�j(�h����P�2�����Z���p��l[����7�rr�����|�_
DK �ulGnvi�6�n����-! �k՟[�Z�f�Ml+a��yk__s~_W�z�aѳ �b+z�b�2�v��8�q��X�J��RY}�@��(�tM�W�f��ǈ�y�s����+��3R�Ez5M��&O��1���N�<A���Wd�ߐSWg�1
���"*��9^wIL�Q�r-h`�ΦX]�4�ևr�/��80	�5�m��#"l�3�:��Jm������rk�7����K<�2'p�p��d�?�x�����1�L�o����Ě���V<Z�,q��哚[�^$%�)r�}HK�8D�����d%�fךo�)�\1_�b�b���|QJ�M�2��c�D�5���#눜�C|�_���D��KP-��s �;��R.�����"�¬mA}L,�`��~:F��v���	)lSC�Pf����@�4�M&�*�0`M�#�j��VKmFD�\��&���Md�.�\9J��w" �H�	A.����{�
��ûݟ�\�@t�U� �����2���0�d㑠R�
T!d��K���T��`X[����������s��-_���~YN�o*�c�M��1/$,s�.�V��
a�	�r����q��w�w*�!��J0���J`<y��yZm��yt���p������~�/p����Fނ�^�-�������#[�_]^�"P����9�1�2cU���'�P+Ă�n|�	f��ð��\|�I\��fTb��W��Th�0!���&V.���%��s?!�|~��c�o����n�Z����GW�DI�=�	r}�S$�1���u���۰
d��6|���.��p#�V5�e@�t�e��	�1�74i������4�*�����j�z/�	�E>uS�`�,G���@v((�Bm��j�V_&(��$
;灁Rzg��A�� ���ޯ�>���Ѕf���GA�MÅ�[cZ�4�7���2�	.�>խ����k>�;�(IS��ǭ3&��ƥ�c�[���lGT�8�'�`�03@�W��H�,�	���:��B���_	�*�7��D�{�!<��]�|3����zs_�h��K=���<��A��Ԍ�@*�Zh\�k�˥��d��6�q;ף�y�
�_^�_GHݣ���'(����_~���h_`�E0;]I���t��Z�ܾ�W��ꄜ�T����Sz��<���n30�O�D��J�^�\��j��߶����NS�����[�by0n����0���Q�T��w�%;j�B�; C�'6�el,S��eⵙ>a����A\7F].��eU���u�#�!Qv�h��?; �� ��8�q�F姌�5�Փ�����H!Q��*!NU�	W��o�y|5�
�KE���:4[��d8d�g�<�'ѓ�� SX�8��ƣ�Q��8���~�&�H3T�`�7�f%/QB��b�<u���3]�S����r����N��x��I���	��Z��7�4��� S(���3d���#����FKp��,�9e5��N'�24���Jӳ�`��W7�`ɟ�
���4`IJ���J��ܙ]jﶁeN��Kϴ5�s()�gv	�����S�%al��7��
�wf��	�_��|�p)�f��:&��V��Wb`���5vwR�S�����=�E*jK,J��ȶ����#-"ۿm���u �B&<�})�t��
����aƦ����D���$�ݡ��W�8*�2�U��Y^�&��	�T�����a�X��s\z���C���BU���@��m���>y�� S��^�5����f�g������i��ڜ��iʧ��q�W����R��!�k>�PM{��D�E7��4��=�KtP����6X�\����D+�b��2x{���쭀#F����K�;�!ǺcU�E��y�s��C(ח�6b`��D��S�CF�4tL��n�;l��Ja��gQ��z���ι^3C��eZ����^�_��ܢr��$,K�kT�~����^�v��1��c¡�f��uı�GfW��Ԍ&,�5���-��?�`÷�2�G��z�ߗ��K^�Wc�����R�W�F�H�n��
.���b��\��:'�aq �1��+C;S�%1Z_���
�?w鎏���t�:2��ao*�I�NM���')��0
�|���� w�cR,�{ �1���<o�Kc��68��������2"t�\�V�K���&��O,��z��K�t�oMWR�ۖ�'�Ϳ�y�=+�OJ�;�5*��9��(���C46X�榹�;K��A�Gb8�k�x��RP��}D�7�]jӔ�m�\�tb��D@��,н�?��aw1ۃY�/��	� y�JE�Z�)�����x)���='�27�^ES֚��M�,Z7��c}�@����I�~��5��;4V�W�Ҝk�Ct�Y��=+�>��=��hոP�'�B�9`�&#ʹ%6b�Iu@�v,�5P��`�n����%Y�]���:��sYu��{	+ =Rl>{}�zAX�Q�3�(R�m���?~��B�zc���>`KFY����J�4���t�j�l=��9��ɒ�-���,����Lp��/n��2�����P�T��*�:V�Z�i~��H��,(��:5FTzYWx�|����G��N��y�I.j��A�h����E�.�6ta��唏�$i�q<o�1��O�b�F=��u������w���{@m�n����`ϯj����s���J���8��q�m��,Y��j��5���2�Q/@��& ��
���#���6[P6�4�e��.�*7�*9\$��������J���n����/AzpaE�7e���
M�D�X�t��Mл��B��ȋ��4Ё��Z2�n��$#�/�����C�p_Ρ"7�EF"JhD�ơ�"V�6��~!�S��&.�5uC�VN����+��:ّ(���$W��uz�S��g��=�p�
<1}�E�I���Ŋ��/ڵ5�	X��L�qTN��#���Q��v�m&�Q��"Y�_iR��;p���&�`F���E��P�AĪ�a��vZ^�s#�>/��!��i<��M¸�Z�23���`�I:��_�Q�S;�?͂#��&�ɹY�=c��Ew$�(J	!"O�`]ܣ���j�k��K��:���A�N����c��D���&4�(@�����[,-	m4w��C�#��4��aq�@��}bd�x2������}�3x5�iq�B��<R_�V�]I*��]�k{3���V6�b�_ؗ����)���G�.Մ?�9o#{���3c���h��d�ȴ��8��GD�bєZ��	��)C|AG7,Zƚ�'��0cC��n��_T��eEC��(S��ӹ�>���a-��眧E:�����8��pѳ�,�Q�14����:�z�|"i�x0b8r�����n��W�g�_���R��ݩ�{�C;�@�A�֧1���/s��G����?�3��a�_8�vQR��O-L��c��"짵�)�j}8���n�l�u_IF�?B���˥yIb{`��w0{�^@�*kK˄�+,Ѧ���?��#5�}
B0dN-�v+Վ���c�#2�Q�|����>�KBU�/=� \��Yd�=���{�x������f�-k�?��"���^�.DIRX�0%ɯ	(�h��z�A8لR[N���1h�}���fE��0/��c(2i���G|_\�Q�R�vb�#T9]�O���K÷=ZHm��tw�����Ze�<��+���f��uj����_�� �Ғ#�[`[��l��j�umW/�Wt:翬�OY	�V\�h?G�����VW��D{���%x�{�a�k��e�Cs��]Bݡ�)�S�o]�AC=1#���0D5�fmTf��	�G��:t��D|���-�(Hw�;���p��)����#��'4�^1	���#u�q�It��{F�*�qƇWD����"�6�E�4	��ѥ+��b������<�[7v�,4@�_��~�;�=���?��m9�`�r�)�d���p7i�ϮF��E1��@nug.�+P6�j��dΒ�g��\=�ޚ�u��l�{�+ȋ51�e�\�H^�'�,D�X?(!�'�`�j��?�	�ݩ�����Z�zd����� E��i��, a�">)m,�Z(���g��H���L����:J$�k��$���~H~n;���a���GGm�16,��HW$�������ȼ�O�
�8&v)����;��t�w�D��WX(ҧF�-c�Z�3y������	��8J�V�薡�Ċ�j�X����h�����v�T, 4�
�p_����l:��VH�s��q�jr
��!�l#�B��,�\�a��ȾG,�i����^�gzZ�k��K�p�i�D�+2��iI�|�8|s��NF�S�f[Vu搜�Ǐ�Ċ�E�0Ȯ�;q�a�ó��k\�|����8���u�Me�VUjM�]��[Jx�͹8^�c� {�
(B�iIew�B�'$O�o)&0�e�k���X	N���Xc
\�1�<g���{,j_j�~��+���κ�Ng��� ��N����x�����-�f%,����	���s|��>�0 a������|A�cL��C*Vm�G��G/7�F�T�H��ܝ~�$^9+�Z<״�RAEB���Fa�d�/��Jna��� Y�Z`����S�����H�|j��נ	
i'vqf=@��������٘@"qX��,�����{�j����Ϙ����~��A=�Dri�Ρ-��'vi a�g�6$
D� a)LM,� ��j���	>���֎��'�!��{�4�f���!5�6;���4Y�r�fv����^�3�9�Y�i�����ٲ����&M�q�"���4�~�cKb�ilӥ4�J��ڔ~���X��4�B��	��0IXD�ٕ�	��f�h�"I}���ެxIa!���X,-Y3Ω�Of`\S®v��lw�K
���V���)�-��Q���!
�J}-�2����A������H���tR�����ڹF$bp��n�іۛ$��+��y���#&<mӑa<N�/nS����g�p�������g
��P����]�
�f߆�X� ɽj�ؗ����D���b�i9b�����5v��o�M�+�_��y~CD4Im�Sъ��q^��2��$�)�&���Fŗ�H���8�]�8wb���Y��H�!NoZ���K�"�?F��.l,���4{�s���-��(�|�pO���6��3BEg� d�����a�<s ��=2�q��;���/#ߞ$Gzd���e�-e+�Z�͖��"��~�o��_��m��5�!}�� ��۞��[�߼�u�s�R�Y�V�qe�����L�ĳ?�is�{�b���X`/�i��߄N���8t�������S�6����Z&�SŬ�u���a��J�?~T,{�W=�8��L`�.%��f}Cn6{"k˕ҾAc�X��<��|�w�wX��,P$�/��MX����LQ��IS��٨�P� �dF�<�ր�>�ݗL%�X������hϓq3|0�{x-�e�״i�>��F��v�{����֐�,u/pi��8�bP�z�H?�E
���}�'���>�=� ��ϺZ�[��J���X���!�
 �z����-��ug���6�7`���'�ë֝����ͮlV�C��Wk�Z�1%D�r���"���X��?(̗�D�Y�I%e�����F?�A98��+%X?6�������d�聎��F�%١��y=�����Y,��i���Y_F����=vf8�6���w�l��z9�=��XQ#�Ѭ]y�y�$&���ر4	諍9���ĭ�uCv*٬+Y�h�����p��ٺQ��Fߐ�l�89b��5F��o_:�	:�]�f�R]&R�	T���N�-��^rͻ1U�]�x-!~�Ͼӝ��;�?�*�*!�j�6� �;��n�%��͒�JA_
6 i�H )H�d�)���Va�[�M��uŪ?� ���=�\,j{ʕ�n�����U�s�f��mJ�&FO�qE��]��`�`���}>~��߼�V`)[��L�F���-h<�x�Y*����"S��-6SG����*�s�q��{����i����<b��?�^�������I��V��7Dƥ������'��ܪ�[�W���XUU��C�D/�(�<qԏɖ�yuf�4J�ac���z����ܖU�b��a��-C!������6�$�D����,�'����r�!G����%x��J�a��x�y�=������}�{���t@�	.4�}�>���6�Q��={03=�w5�q*I,�`Fټ��׿�|��k���y���zָoc����;K���B�j�o�j\�N�����k�@�y��:W	���؃^)yŎ�HCo� sV^�bR�/G<ñ�85c��E���N�<���u�7!�a�x��ߙӑ;�	� <2�`�C*2���.��8��U����U2�]�X4&[�_j���٭79XAY\�CQ�;�u[���^g{�:&�<��;9?� ��̷��s1)�ڶ�����i�?۵.!cu���(�V�=����s�7 (�8f����"
D�x̟Vߚ6.�;������w�0f��gv���wP}:����KT�|`�徳���^����pRWQ�/���߿��u ��`�R@�[��6����)�b1	�g-l��_,�K��A�>�NIfn6:�eg o�d����5B�-p����1�
xF�'�4�e�V%?��V^0۰/��u��?Urrf�!X.E"5;��|��_]��:�yݼ�,�I��yBT	���b��ʶI�n��4c`�z���m
ڨ5l�Ȓ��W�������R��{��}o�8�2x�)�k�	mY)#�.�oO0$����Ө���l
�:���]�,��뺬�D�C�:��5�֎xk_bdu�%+v�?���A8n ���Agk<Ԇ.��k�kJ��Z���=�]N)���� %͚��@D~����_*��(�9��V+j=�)XU<��"p^\��^��J�V���N�$��k�V	b5���Զ���o�m���^=���9��D�1�r_߁4m������&r��_�i�qeq�s{>��J�xv��y:�ZXC2r���i�6�4-�iH:_����u��<]`��
���G|�%�-}����th��ጴ�@�k#O�b������`�m>G�wpz�s0v!S�>���q���4���E
-X� ��KB-��dcoO������{S/�$�m+:%�uo"�j]z��;a	��~̷���I�
ș�� `G1����C�VA�I��F���I+�����T�bU���&�����	g��GFm0�o�3�x�� �(��o��wP2x[x7�b�2]����m�6I��-`z�f7��'Sz�t�,�%*��Nd��s�$%��2�e��M�u�h�!,/���^M�O�s�R�X���z/�F��{��p�(!|a�Lxq�f�'\o�(�=��<���p�P��U��s���b��7c����x	#ЯRjpz/�(�8:Ъ�d� m2�[؀��k�����9V�&�N�3��|��}��$PW~���$c��� ��Y+#!z��t���Ex��y>�5y��̓qN�8��ln���QpS��4z\�9-%_X}�-^��T�HJ��<��j�~o1c[�l �n�� �j�4zi��YYnu?l��F���x=�4����ZD�[B�D���I����ʯ=�s}z�l�I��o�@�D���x�lgW+�Ҷt��˖ǌ� BEl��g�4Mn�"w' fT1���_�䦠�[T�s�A|��S+>r`��'�n6Ͼ\�P���{�]�>��QF��Lj�1���$��@"�]��|��|��v�ك����T �������18���#5���M�v'xR<��L����s0��c�rV�<K��ؑE�փoC��o���Nگj���Oa��IW���������t`���W�@Z�J����]J[��c��j�9��j��J9��Xє�D����zŻ�?��q|�q�ܩ܄[�dh��$i@\���.'C�h���[=���oɬEz3��Pm�,��S�@�N�l�ep��XZ� �i�Ft�{�l~eΐ�����~�:�-�i�0�#�6�˲@���8��
B�_��C]��!B}�����]Au�w�-��m.!d��L��QK�6X�~|)y��x��/B~��w�b�N�
���2�G��L�6=�%�J���s/o��]�Vu ��db������(2��dX]�K,��a��Q%�|n0J&9���=^�p�#��&�k�5=Pg'3ˢ0�Ï�]����yv,])�8y�ҷ��z͌)��=�ޥ����z�����c��f!��)�K59^n��v
��7N��<�l�y]y���֒�	��Y�s��A��v��F�X�(�e(�����z�Յ7(,e�&m���-�t�N�AA 	崿�[[���K� 1�G�n<s����p�߷0���}\2�+������'t�{#�]W�`q��*��uq3&��xY|�lt��./�!Ё2X!����G����ޑ��� ��Ld=�ȥ3�H�˝ڰn�. )��]t��3���JZ-�֍�c��>L��P���G55aDC*A3ĕ����:�.
���F1>���t�� 9K�j��&O����= �T��LA+؅d��o:�n�������C���l�dws�g�.�R_�����B)R��Z.���=B��Wz��Ґ���_�V���w�rw�� �rw��IvTG���6O'�֛�\��z��m8���f��+5`�B�~���[��-~�k̈́��4����V�ώg�R�2ʚ����<���S4�~+�E��-�h�m��:沸s�ڔ*j�~2D�/��id`�Ql���C�)3��[���8s [t��~(�]�T����Z�٣W��S}��X�3b��?��?�k�t��D�Μ����grã�_�N�A�I�ȶJ�������\>C��}�����f�^�Ix��n/����߇�"���J���5�� �h8���V[ǝ`n���O�#>t����f?���� ��Gy��a�Ea@I4>�J�P�D�R�ӿ�Ťc��8М�p�x�	�8��N�
�I�
�xs��`��Ip{V����qc(绢���ƿ�i�ge_^��MM��'������i��u��&/G׫��CX�e����lH���y��S�	�xG�oC� ��6\!��;ɯ>��^o���zvD�V���������I�حf�*t��� /#���Ӭ"�e,	m*9�Uy9]ߩ�&־@��Ͻ�o&YIdu��<�+֞����o�3d6��}%�}q���McE��}W'�M<�*IXnFѣ�,��9q���xF��c7��5���	��K����V��I��!h?�����>���Ab��TF�Y�8�>���������B�m�ߙ�x��e(����$2ѝ��]d����Ћ{B�C� ��FI�lG\|鞌s5��ǲ3�J_h�t����M��ުҵ��gN���	�Q���m����p��ӽ�_8�O�����"xu�M�}��F�f�a��i�����E"�t�Ȼ��eT���e�E��\>RP�0_1�l<l�z��Q	����Aq���2�x���d�:OQQ���e�3�w c�m�^ߝ��%O΢���+��8��V�������/�"���2�a��)N���g��#L{a�E&O��_I���f�dSR���<���h41N:��R{��=�K�W<4��V��%Ug:6�{��	m���ԌH'B��L����m��L�>t��*tp���_�Ԥ旑ZG�Ծ��f+y"@C;��e��(��ҟ�	��g˔��Pf֬W�#��a�6���-�"�V�D�J�<��H6pލ?�@'�Sv�!�Ek��.٦x���!��Z��eB��uU��p*�����uG�����4��y^[%!��<U��|x�U��l(�EZ�"lb[�lCJ�{���ۯC��=��4��egsRbRi���n���L⠮+D��x�j�����L<zVسY�ǈX�!k8�8��z%���*�2�h���`S��vI�^"��BMUq��hA�@�ֿ8�a5��ا��Z����|�c;�{��fb~8�BAGyg��D�kF�7��Ni��\&!蝬��J%�v�%��`����?��dn���d��nm��lM�`�����qң:l ��@?�4���]�&�f�����L�Ryi���A)��;j��?�Z��?������ o��=hn��	7��e���� $ҿ�k����j���	z�ꩩ�EC�}��|�
��! cd��M��ݼ��1�<ڼ�n�K>!H����}�§7�M�%mo�~z"`|]�g5z�X1���pg���6�AJ>�I�>��g�ݬb�����{������C4��ʻl���p���59��~��w�0������##��S�O��)�Vuj�WH��m�S��&dҳ�yuKN�ù)=^�`�|�<Z�R��	7�#A"�9}�aq�ֽZ���"������= D���M�����x�@7�q�ip���@���E�F 9�ݺi�LZ����0t@\taYM�Ҏ��~��l(�,�ϳ�d��W�������fٛ��'^��9� �^��PXm�.�b������?��k�6������6���VI'�b
�.�'�N��o4��j�~9��ORr~���vls��m�5L��^�T�i�5���\	<^;�8����q�ѡ��m�yboo.������'Mp�J9	�m��%�k�l�?R�cC�qyVl
�:F�<7R���)�_�ŴF�ɂ���"�2@v"Y9h�e#C��Q�{6'���Br<D��h�&e|�;�t��I��/���4���in��\�3�����O�OF���h�|#��>E�� �D�k94/�[l'M��T�$7+��U�x�&����7<�d�J������#*Ah�`Te"���fT�%�Բ@u[r-�K]�*��y;a�j*��,d���Яk�[x��z^���/]�� ����t�7>x�"�V1!�g��L>N��pIU��m�z���R4�w�X�U��Y�]�YD�%ps����F�6�u�3����sH�૥5/�`��|(Y�$�:v
ِ�ry�n'����H�A��"P�D18u�A=!kCnf�(S#Ǡ���f����[>'w�����=����<6�`�s�����|��A�*$�W=~%gDb��uoy;:�z;���0�	�R��z��a^3�ڧa�}V���vǏ��St[g1q��	�T!�^i�B�<)��G���0��z��2c �+5��xy��K�8��I��ڹE싾q�8��2H����9���nC����� �턞���C`+�A�W����x �T;�R�8�����?ǔx�_0���͸�U�cDб��%y�`�ӱ\��Aݳ�[חX����P�7dR�����F�ϊV�q]��`p��C}��VAg@ʅZ���ؔ�h��7
1�|�C ��&L��i�T�A׺E�0�ضq�/��O\��)�.t���Gx�Ժ�^.��5մ&�v��l=�!<�zQ��b�w��:7o��:�ώ�*_|�j�:=�ù�:��0#�9;R\��i,0�#4s����D����t�r�>��V]��1�&H82�Z�{$Y�8�]��pB�"�v���H�c�x&\�	h�^\��WY�>*m��efA���k��a�x����o[�h��� �Z� F�Yy�����$bz�dz@}j�-�����߬Ճ�ԺEh&�`7Сa܎I�,IF�D�F�4 �K3�����\+�O�u@�����6�HM,�U8J�(����0mU�|�m��6��Q����K�w�-�خ��j��QfNS¤v�zg�#�����Z�J/���t�61ݣۄ�P�1}HU2N���1O����u ��FΑ,��ğ	z�I
/���?�Yc���u�4+c!<Mx5�\���`��w^,�q��Ozx��JZ�}p�/l�gm�}]� ����D21��T��>8�� ˂���#�8���bu�Y�<��i��?%lF��SI=b+}�Ԣ!��]��D�-��������M�9��-�Q��	����,^�#��A��>�:�|�R�<m�/��D�� !�����aL�@
ͮ-]a~�������p,t�Ӈ݉���_^K�;Ԩ���%Z�{0���K�4���5�&�w-��)E��Π��Z!�9?L����1<��x�4y�-�kD'0���5l������zΈ��V3������s�#�e��#�*�K�hY*erbw��fg>��	ڭ�41�l��K-*|T^,]dv8��u��oEz�eɟ��LB@(]j�U4@mYp�ȟiӮ-$���3ǈ�@ X�~~N� �(JT��,�Z�� \��#�cqp5�Go�g���#?0����o%�=UM �Vݡ;��ńѐ����V����7j�K�3���yg���CB��"H�[^@!vL��\�oBW���������E\�Uw�ϸ�i� ��<|>�����b�&��-�2���?����>�ھF�7�r�l��/��`@2xv�A���\}�-u�>�`p���E�C���"�#����Pqy�S�4�*�S�������{�� ��aNv1\�A�`բK "~x?yb��<Yl��&�ن��ǋN	��v��|�a���(PK� ���6�����
s�������1��F����m�%�O�"u�����R���cK � {��؜U�ëo31z&�Z|�͕7����Z��%V�З�w���&�M�΀��S�rO�X������x��b�'�q���B/���ߛV��Id��&D��X�$'��k��d[/�d����)l#��d7��Mg:eh�?��f�?�5��a���	,gYЮ-�#:Ҙ�&*ӱ��Bݰ�K�`��}��y&u/���4�q����Vp��,aD��x~��C�JC�9�������R�g�@'�a@��4��xn>�N������Ʒ�P�\�ǉ@s�`>�R�t�Cz}�0�+���k�^�)��V>�U||� z�ώ �$����˯pP�q�ǚ�4s@m������6N|�d�$)�m��ȹa�/o�R�N,���	�'.u�e.٘<:xD�=۟�(��b�����T�� 0c�������z��HԶ����?)ͫ%P� "�Ae��4��|�.ci~uM��Ag h��߬�t�����.Cj�O\���_��m���_̞6�HD<�|a�n�5��%�BF*}x&��[��	�$�?����e����&�ߺ�~�?�F=-HQ�|��Z���۰�H�ZOa��5���L��t���$�	�a&-Ғ�n���a�����J�|\Q�%�=�H`�AC���YGD?
$�:j0JYk;[C=`�=\fl�¤�Uv�i���?��1�J�����C���FZ]�?�2
��~�	���f,΃�+�	�t�~��tr
�"���u1�z����]��!�x�t�d��F�=p���h�g��`���ߣ�	�-w����L�H=5��q�ir��Yҍ�<5'����=�dq���Hp���vuD1���-|�ّ���N �O�.���%�3~r���S��kj�Q�u�<I�Q���uALx1"+�5�Y���I�	��/���ʍ~h�����ڭr�d���)\3-��]#p#I�QVY�S<?i������=�^�P:�:����+4�G�~�vߘ[�m C�<���:"'"�G�3�P���.�1_l;sy�`w��C�e�ٶ�Scta�ѦD�����@-�|)��y�Dn���P���ǳ�ǽG`77�ڠ�� ��x��TVՖ�pp44��&n�UeCaJ<��aW�d�=�����ٙ�5�%��4K4K��*�e�k4��Se����2��1%�!��ds�jt[�Ra���	v��Xf\�r��VT�-"���Q��\�̺����s{:{?F҂�Q�A��+w�-O�����rdf��2����"�y���lGD9+ �1��i��V���jS,U|vag�U�g������m�x�q���4'XWJ���d��k��2�W�z2�đ�&-���z,��,�	ސ@sˈ�fN����1z�̩l��X3G����j{>̚p/�i�"�ۧ�������)�����u"��4d��q��n/���."=��7��Y�����s{�����P1�>��+�3N1<K^Y.��<�/�@?���e��Ƶ:�o��$��^�~�H	u�3J�}2�_�CFi�X��V�/0�ўXp5f
A��n��DC���4ź�!Ȍ��\�.��nć��qg�l�+�:"�cĊ��?;���I�B,��_�����Rl�,�o�=�SSڙ����j��Щv�8�;�X�m�1�o)"�J�<��֋��!Zd��G�gOY�m���gS��)���=j�ŕYBC��:ԯ%� ���Q�8���Y
ɾ6V�D y�o/m�$Õ�_�v x��h�_~-�"Cm[�Vd����@Ԋ��^�x�}�ʢ�J�t�r�$�''�.����$��ƪj�����T.���M�����hK���W·�27pa���Iǣ�� &qJB��o�����7'E�\϶��8sʔ�LC�A�[��ART�?��m��n
ڌ�u�6�sͤ����B�|�`j�v��%{��0YD�G� �T;�	�!Q�E n���8��������R8L);��E<NA	5s����C\�m=<���b&����d8~W؀�D
)����@��[���%��p���nR٦I�K�}��k1�e8��ԝX�jSk�Q&n�Yә�0A�1i8ܪ�52�j���v��T��;���^�_՚�{���\���[�<��.y�,k�0���]J5>C���/��A>c��	�@��~Rf=g��Mo�W~�pl�j�гC�qZfKf��k&����)�3�دŤ�6ؾ'#�T����CE���c��DF��9��M9�F�Z��5mFE��R���h���6D� ٗPNywW��l<O�fJ>#�����%�j�5Y/�_�7cN1�U��<3�C���K��,H;�;[F�h�ΐO\^~ �^�`#���C�&w��
(�}�@��>�P������r�HY��D3� x�+o�t�1����NQr���'�t!�Q�܍�Ʈn�qd��jTAZı��:��~�D3?9��(�⸥
�l��
v����`
�����*+K.�����G���~W�VruɅz�!�c]���Om���j���> 9����88V��)��'�� �L��$𦾞����xXQ��u��G��y_O��q������&�E��o��"51�&��0�O��+̑���2�2�?��7�_�$�$o��F���k8\��Z��D�M�� ���,|���IA-m��{�&���AHb0� �6��P��Y���G��g��o1����,G� �����>��✌G����Z�'�]H�B&��k�xa�Kѥͬ�u�7J�4�n�k#1�!�@+�BF�Z'�c��7r�����.��h�7�mW�WY�(W�?�:�t�L��S��ՙ8�x���UGL����'r4�0�e�o�#</E$v)y��N)Y�!FX�@��.s�� �1��h�cXU�7����<G�$��I1�
�l��t0�����v��NP�*��H�0Gc�ˡp}����=J��s���-����:b��-I���&���4MC��Ӹ�]�Ň��,�)�W;L2�-R�!0lLt� ����_\�T��v���)F<)%�o����D�T��Z�h�`��,CM��Y��<n51©r61������h���Ck�Crv2�V���#�����ơ�Ƚ�>���`��W���ɷ�*	d���Q�鑂�s�v�@.�A %�kC�O�܅Lrxe����	�ʦ	I��.�8�׼}��b�9L�#��c�{���J������O���hx�{�<ӷl�tg�0R�D������x�o�"֧�_�&}�g+���I�"���&�H���Nw8`������p D��*D-������Po����.eH�/l|c�˞c  A�b)y>����^���Q"�|��5���Rg�_s�S��y�CϠ-���o���+�8�.�{�NMmBV;[u���IAn	�^	��|Vn*r�U�2��;G��+��NJ��	2[�p8�w�c�������)����
9]���"Q
�Ih������ٹ�S�S�ì��U������^\�}�'��xmRh��Wl�38���r�(S�')� ��'��h���ݴP��d��~#��0v�Λ�8��c�#Q� b�� ��v�D�{j-T�若�2im�; Z1�a�z��czj�=�AX�� �3�{+2۫.�b���D_����Y�R���,����[9�Z���gIzN�3y&?���2��=�O�s�s$B��x��b�>�yhF��Q�çb����h~�2���	�������1���H��jpY���Q���I�?9���G9�j�,*ʒ|6T%��-R�`����`�"�>�{��A�5���v�ɰ�8&��I��n��샂ݚ���W8�}��2N&y9)��z�����$����U����v1�)���ܴ��y�������I; D-�0K+�'OEE%��m5^�xUi�0+�ޖ�N��?�~���_j�`~��i�x~`�Qo$6���8w�IwRM4�S��7@'�"�*)���$��
*�}�f�������3���?�F�� ��˧�a��b_L�F��9w�7�ai��wI� ��s�u�zir=�>�s�Jv���;�͖�y;n$��$}���G�<%�v���0w-�Co�c8�6+�j���O�%W9P}߯ν��u����&Y[m<����<���_�x��n���r�d:\���+G<�G�p�B��}�Å�MtݵU������dʽ�U�7�u��i���C�nIJͬ��+���'�ˇ�^���}�쏋T`|�� n><�;�	�r���=�-���BrY�%�"q.Q��0ܿ~��!��`Q}���|^���JY $��k���P�H@�D���E�qZ������:7��B�)L6[�����r�06k&����������o5�~>�EB�am��ݟ���\Ѥ�-t�4�b�(�Må������F���zd?��4���W \Ҭ5?�X�t��-Dg3<��T�� �j� �m��|�ȼo<H����8�0���q����L qc����&@j���V�8�sI@$�?�4���I�� ��<m��\��xd�������c��V�8�}�e�H8�D�e�[���?����	�0���,$K)��Bg%�~�/@c{XL�Y<۸�8V`
<�^�.��7�}j�CY�g�:�l��yt8 |��!�r��QR�
�<5�>S�cRtH�
b?��5L�B`BE�j�^YX��u�
;xs�`���i�t��Q�X��؃@�R�IZ�mf�(�_;u�rч^�Q�S������,�3G�fH`]t����<M��y��L|�}(雘����'އ0�/!l�KG��墌��I+��ڙ�질r�8��Ѵ�*�+q��ʝ�W']Ar�W+}n[{`�m��s
�zGgJN�W2�����89^A�l���|�V��+��SQ!�%�	ǂ��I��f�6e�{��ŅV�а��q�ò��8&5�S�a��0����|lvh]��lk�n��ݨ�@:�lhC��/�rT��GS�Y�I���Csņ�?],�F;�,�)&^=3'���1/�֯��s��WIF�qj7rxyx����,T�|�I�������������ڐ
uh(^���qk7+j�MS׽M�;Pe�6���Q�|iG�<��v�!>���DJw�7QD�,��aT�E���-z�_Q%�8]g�(�k��c���"7"n�<M���;����%�o@�A����I�'!�i�겈\��7���`d��k���q�q�!�L���w�X��F �E�<�@0V-$�� ˘V-֪���8�݋Tl��'�
Ҩ�e2�x������}��k3������^`��p�YA1���ʸW��`�� ]Ŀ��O�):]q��[��� !�i�fE����'i�n���
�g�.�,�&Z"Nێ�|a���%�T��T��&�<u�ɮ�0��N���O��:"��8�\�B�-�\ �*��*C��Mb{��-�ֆ���=a�ڶ>�u$č;�U~~�K�)h�_���i�VxP�t���
�΅�lۈ�4��:�hn�:,;�>��qJRTLVb�R�[dWhN�*A6mץROK��5�m�t-��j�.<�c�v�g�X����|S^��~1�SW�)�\G'�䉀~'�F�rmA���1;WgB!�v�'��(�deMԫ4o!�A�C;bX&5�	�5]O���ꨆ��
���(_�l��qt�uQ�	M�Gr؈(0�~�*��_δB���VB�"�P����uBGUŵU]�J"�0no�᪦$�X��,� �w@&j��D�+���Ww?}��AҰ����+g�"?�]φ�g"�X����Z�ܻ�!!I�̄���ѽ�'�����ց�T��b��xs��o�l���;���'R��M�$�R��X�4p�B�#F��1�ME܈��sY��3=76��$�Ak��J��	R�/��\�����7rcT�V=��0��-AWةk)#�1����x�#5����_�t��B��YK�<���0�,@{y#'��6���"�vH:V��&.���������W�Vw,^,��:mg&��m*�Z��Q�C?~�2嘎`to���j-[ 2���E�\z��HxސNu��/���QanX.���o��Ð������ʝgx�51���~���=�D/W�~z�7��Q!���`���P|��6�z8���t�(�94�\Xb3��˯]�{��ϼ�nt��3̈́���	���pX��k%��M��p��%r�\Z�+��u��Ko��2�(����\�5P~8����[/9��5�,m%.ꥬ'/uU�z����2Ƀ�U����4�����<D��-�^�P���h��՗L,�����ana*�����k�!.�F��7���/||$u_6Y;���������p��z[k�Gdd ۧ��6�G�n�*�5E�А�ƫ���؎��/��\��?�9�B�ցj���\��R"�Q���4���5}�`.�\X/?J`�
 �`v�#d���Z ~"*j��f��P��R�� W_�aޑJ��H.ݿ�]k��
��}�M?
ͪ�O=pg�l����˿Wq͖�!T�= xi#1V�M�)�=��8��FH�-<�k�f��� ����B�nh�s�	�~L�[걜P�d�h��&J�X��6}��6~�@�PW��M����+�x��x���J��_PE��.����-V��8����J*�I�ӕ
C�����bu!R�;��g�QWC�p�lkS}&�$�mW�I]�|꼾f�
F�<�J��V|�W���}zޏ�87��١�Z�U)����+��Ok;������zJ��N�ٗ;0�`iPj�I��^���K�(��߱�}[�p�G c�6�(.Sû�g���gX�G=V�탰�� t�����#�[�a��m��� �D�y�l�W��)�/#U,|��\u�����0k�g'�!+������d�&������$A�^+����V�\o�\k(���HwFe���6��	T��n�5�ET�Ȓ�w�2��|��̼w$_vق�;�6�����3�����s���#��;��y1)���8�x�]��iTUmd�V�2�<�֡W�3���P �`��Z��37�F��l;z�
�5?��\ۛvS]�n-�|V�_��5=��� ��!�y�7Blp@J���y�'�]a�A�ա�n��Sfa'(j����֣��*&(���`����u���b��y{�Z{�+[	��F;�LT5%g��m��9�Cł��/�Ģ��LCs$C�sTpݒ�a�M�b0Z�#N��K���J=� �Ž)�V(�� �o�� ��I�y$�	�J�'1x;���	�;��V �(8r,�ɫ����9K5����3��g
G
g���������g;�x=�����>�٫9�=����|ʚ�:E��#!M����gr
�l�UN\[>�_�'��l*(��G q�� �}`}��&~�,Фu�:8��7�S٭��ڎ�	��j*4���a[ Tx�AhR�|.P-����	���GW=��m�޾�BB[ߛU�Q9��B��tg�>� ��"l�M���)7� �����{:��ꕒ��Ce�(��:��b_|�q>C�|.T0�^V.(@�� �S6��C\�?DK���K�ҩ�CO��?�Y��|?N�K��z���,P�agBI�MM�����_�w���`�E�7�]�+����� �q��'��L��J�V�;���7���r��`�=�u+���\�54CK�%s4o�c
E*����Q�#b�cϛ��>s�/����ϣ��6��pB�W�@C'^,t���M��I�F,�a�иIS�E6iϛF�Ȏ|βu��Z\y�E���ؖ�UqN�xU������ݴl�O�r7�ɖ�{-���{CD4X��;j<J\�-�z"��r�볯�M�'�y�^b�V·N�Dc�W 31Q��^E�]H�4��NEʊ��1M�7`���$1�:���	���
<��\���.|�z�@�(&kx��(�ss�ф�:Ā{s8�g�\>)��e�
���֯"j�\֥��)�����ƿ����tI���V�b]�-�CLF6��sNF=�y���`"�*�sZu�:�(+������2��zr��T�ףd���睞Q�0�׻e
��R�b�ūka>/P	��3[��E��+3�ME^�\����������JCKI����x�":t%	�� �2���9��U*+�A7ڜ$P�ZC�n}��*�M� �[_��joN)$a����B��U�=k�O���#i�@��u����2ی�f�7���a&�l�E���d_v�k���4����N�@"���;�bw`Ĳ8�� !R����)nD�v��yq+�!;�| �M�����88
����$����^d^Vdmk�i��!�B�,�
H�tDU�%�\�:xv'%�b|�^F�����w�O�c�`F`��Ɩ�ґ�(��]�bx�ݼ8FC2�5|�U�kߋ�Jꎸ��������9�� ��hP������A-b2d�)9��~Ȣ*0�<�D}\��Q�(��w:��]�4�p���#����)�3��ġ�$����=T��������ymȈqh����w�x��ɕ]I �n��	�Q���ЫN�Gd�/�#��ʆ�"fW��<~���T^A"��@O�	�"���i�c�0/�^���2�.,�M���ux��|ru!�n1�4{�[��(1�L�(F�|� &�b�$]���'L��	_��v %[;B�7��Tyټ/�m�Iuhe�btn��>9���X�%����Q�DKZ���0�;�1^�aagfX�h�����D������G��
K�#����LX��v�Wܹ�2|��9�F����ݙnm@s.+�a�$��C&�}�B���ZG�@?�]b���|X�XZ#|usH�C{�t}�9|k9��6]T�Ex�^>j���D[I��[����h:�d���l:��{�T���˓��=]�2K�����P����%�2��>���� ��Tt;d�L�Y�C��.��� ���!��j�9��\ة|�j�Oz��&:ik;��m�2�HE�O,�2W��ql}�Z%yt_�aWv��廙%��ݔ�R�Q	�U)m��Ѕ�Ŝ�EN�|Gm�N)~��HX��y-/\��;��\��
�	v ���������2{rb�-ֳ;Q��vg�0��&�w/w=}������u�˹o��6����Ȕ¥��/|�w�g�^��	z�=��;V��o�{Yfx� ���| �D�LUK��)�>�z������:-F�
N�Fi�/�ꍥ�тwǒ�ݢ8��.�'����'!�%W+讔K`���-)� X�
�	�G_A�e�Γ�{�>t%��������fc�J>�?�J�$BzSިI��M��C2����wx�9�9��0<|��#��ۖ�pn�i��X4kW'�o�ϊ�9�2.��2sn�
����}v�U�	�͚�̝�q�sw�D�����FG������R��>�޲Kg0A��$�&���(6������Q��>�Y�Gt=��s�͆�~QQD�6FM�l�u��O8oZ�p�C�1�b��ᵭ��ԿeSG �@l%��1����dwD�T"!\��^�>T��vR<Ȋ��\��npn1[1�)�,�u[1�g�ÄxYUkvC��υ�s6��{ y��Qp#3�ÐO[�Ċ�D��(��%@�q���Q$O_�� e��{-�z+."���h��Ȍk���6�/��f}p�
�;��%���(���#�e'���)U@T5��`���*!!�����0od��xC`���MO��@1{��v;F���{Qi��%h���Y�9i�`s*^�����d$y��G���|?A�	K>��MC�9Q�胣Yg"W��ϩg1�����p��a�殮B�1��D�N�д%�N@��I�*ّ�ҳ���2����%�:�=�܃,��if}^�4A<�~$5*Ӡ�/�9��&
�!,�%��<2ʵ*>����9Dt���. ��3,�o�J	��=V�����j3��M���T�1�q���3��	��x���k�E�s�MJ�8�翦�UF�29�#�6�`����y�6��d���Zvk�x��_�|$��:zf��tH%�>�E��TA�4{s�تoL��D4A���Pi��ď�}��� x>D��G#�_툿�JђV���&�HMI
Ub�����H�!5p�3����Lt<�<��~�U�P�T�i���wK��3��37f���WMkGcz{�1�xej�d�+��[7(�@5/ �}p�Q���h,��y�*jy�<���Q�b�r�����^n]	�������U�����ɩ�Ξ�eU��W+���h��6��	Ǭb>&Q�����qI��~A�LcB3=��T�	X+ĞWI�^��ȵ��v�ԥ#z�X�qÞl1��DNJ�V�/�>�����fp�b&95�E�,�1I�Y�����3p�ۄ�BҼ����P�]i/*� *Э�н���u_�0�������!��6	�Q�aٓE%����J�.[��ZL�cP�q&��k�P_����Y��f�h�j�K��!e�y��6��N�c�)�5�C�{�!G�FqF 3#�jv�o�]���(���NQ�,&�1g��L���_��~\�姩�|ةny�s� ����5�{���K�Ń�;�8�����b6��,0��kKC���+ۤw�~���W�pQ�k������8e�d=���ߵs����]�B ?��]�j@sN�A��L�\��fUwU���7ľ6)�<����[�θ�����1�k����^�x����q�yH�%�a����0A�3�l%�Y��nW���m��'@����������l����TC���F�$�e������ۙܓ�{�3��[yk�u))��q�ի�Q�RQd�پ"[��'���~�a+���O4���a�FXX7�W�rPG�KI�\N�PXv�>�������e}�����_)H�/����a%[�ϣ}8�S�&��S�2o�l����Q屮��gŇ��0$�ҡ<�:Ze4�
���iWZ�r�hd�`�aM3����FEwU���@�T �D�Tl�%�S���&f~�$�L��Ě�V�T��0Ђ)b�ٿPZ�B؛؞	K2�����eX�෍��,+���Fp�e�V|�x5�K,�1N|W�\�������L�ǂ�xݛ�Hڏ�p6���K�� ��|�a�����OFƖ{J�;3[Fx��&剓�7�3�ði�����1)*��qY�욥�$��\�4�J�?��˹L�E%�t�D�fO׈!�46�4�I[� K��E^D�7Ü��+Lر�1��^2�؂h��ֿ�}!Щ~�y�' �����|��4�e�q"ET,�9�(6��C����8۔Z�'6�<�;�'r�����j��ۚ�f�7͛?�g�3�t��䗰K�04�MV5�'���b�������2漊'��=�*�٦��zA�b���e�g��:v�o�z��"�-*�x2~2C�#�4?]x��n;�+ǭnTKΓn�TYݥ��ˉk�B��J��v
���z^<|�[��\�<�X����)Qp�c�s�*d7��@�V��.��Ra��_�h���@ \,�ɜ�Xj"v�y=)�^��S��_��3��o������
��<���URV�WE����ϵ[ m�o�ѕp����my�W�R乻�j����<%L�г�:e���#�xD�˾���ީ��I2�uD���*d!���ْ:�8�4��Q?�x36��ըg��Ɍ���%u���n��Y��]���4�VS,�)�W��-�>�2n�I����,�jNuٰ|��;�~h�f�vmV��+;tQ���s}��b(���`�WO�ޭ��1Z㫋�a�	ku�95m����w�����!C(���z���o��!���-[��y&c\tT�N!,t��T�kd�Ld��㍬@G�qX�gy2;�X�/lҎ%@�^(�0�6����ҐB�L�Eݞ�bz!�
'�d;��mio�bLE��&�U��Ɩ� �"�X+h��v�@.�Z��t���j���dH�h�7� �')�ް���m��r��+W���!*'`:�ĳm@�7��Bci�r.Ap�4֑mNC#���T���'9��\���}YB�-G����N���-��r��|6q
�8���Q]Ȉ�}]-�Z�oe����S ��r�|Am�c�[jT�3*�WJ��#��׊�B˺�\�bm<Ӧ�R�"Kz�R�w��D5+Nf&P�����?�e���
��&���i�/�Y	�[�c�2O+t�BYT�s@���P�Ŷ��",���b��~�´����-,���K$`o�crie:1�����Q�[ l����%�l��,ڶҕ\j_��ǾY�ΓW�0X Xބ������d�+�D�$'�n��F���,�I��P��&գb�Xdk���q�� �y�Rew�#�1��?}sB|��|'t@�@h��#GN
�2�g����I��Qsl�l^u�ښ�Ez��vi&W�!�o4���A�^n.P��g=g*'�-�-�kY $���˨Uvܙ�6I��J��8��������S������.�01�b�pb���,P ���Vb@����taz�|F���q�T9�#�mkN��p��2;u ��.=�}���3�A#Fg�}��X��Bɖ�?�s�+��𠱯�"�D��^�-�<�:C�g�J�N�H\{��v3.G+���h�$��Z��� `��6`��ޢ�3�mrDGý���ZJ�d5�n�¸o��h�+e8�� ��"�/���k���ӝ�5��;:��?81�̷�o�,-�н�x�����f��Zs��w2+�L�f��������H�Bsl$�g��t�	 V���@"dtD�BIa�s��|���hs�IjpB����@H��qW�8��';%Z'qnS�Yx���6��,#2�"�?jFZ�`�(��H��/ӛ�I��q�@/(���\l���j��}b�uL�"YW\�dJ��G�ݩ�Ђ?ְ.'G�_Qtave�������tHG\$�I�"e�������/�����o��H��
�/^��ss��l�I	rJ��*��Sa=�HS�۱��2��Z;�P�x�\�e��85+���s��A������L������-�a:��c��S�`���%*DҲP=���\�۷���ↇ�����E�"d5��˓�gȴ���J�A9�)���ŏU�E	���R3}��q*Wy{Hܕ����mw�A�G	��os��}���ޯ�"�fY]J(���fsP�x[��	��	�<Z�7֟(rI�=Dn�l5 y��e�@�x�)qt��R_+������ħ{���OSYDK��sQ)�ҙ>k�)(��s�CS4(#�'�nw�+	�1�Pp���T!����^ӎ�շ�Dͳ��|�����!Ug��R:-�
h��Y�p<�{�~��B�׮��5�'�������h�w�O�!N%x��X.���Ip��VU��k �ʫ�Q�;�[�h�)��/+Ѩ��+�/��Ui����+f��!�g9ӓA�[�]�}�m̾YQ�|"T�I��ECW]ُKEj֡&���?5�|��Z���2��|����m�x"�D`v�,�G�/�c�uz�S�i���=��RD���x�}w���XK^oM����v��v��q�P]�
1� �9H�2�*�����.���%#Kf�㗘]�A�dxGϯI�w���=��Ŕ-��7s������K�ڳ�"e,�F
��'�������N��8��J�
^;W��C�q@���0=�er��G�+�p�J}TvO���~�� Jlr\��sR��o���R�^�l��!8��tE�l���Jԟ D��\U��`c��Ӯ� �i�)����M
J1�Lg��y.��Ig�[tR1�EY�CI�5w���Hg��Ƌ�Jߠi_�"NRׯR��[��Ͳ�nh���2T"�im<L����LMn�o՘���XY�����8\��Y�8!�g6.�����ssY��Z�3�RP���k��Iuy\���T� �2�]�rl�,)�T�%L�tx'�� 6���z�N8ܩc΀I)F�㎰{N
����T�8�4J��bHK?b0�u���=]	Sk8rl�o��:�H(-t��5�|�M
�hM�>�?���k��s��ұ^�T�av�X����+�B�Z�$����	�W	���ڂ����hw��lF�[F�mݟ�]�[@�n� r[JJZW��!.��L��J����Y�<>�tK��&�1��!��3��#�|��R���@�i���-7�Y��O�S�0|�M��ʛY�!QsY!+�*flq��,��Zb������!�$�-%(<�8B��������D�s�r_c^�Gy���\f��Q)��árQXP���Ί�yZ~�K�:V�i\�5�:w�Pv�Rx^�rֳ���ݐ=mI4)��zT�9˘P�r�q���հ��*��&1=!Ѱ��A��Fv3-����>wçj�%$��Cuf���3���qs��T������d����W0{��u�B��RP�#ylw��g��{�.jM7Քt�?��P8�����O��8G�����e�Wl����@�F�|w=~�j�����uK�G&�� 6��C�����;a�$�\o r!.�'aL��Q�)��5:����xc�[������+q�^�y3�y������.����tad�Wn��`^Ni�x[��{V؛�+�f��ƣ<a _q��*o#���@���l�xVE�*�t��]k��'$@�������A�q�4q�J�������x|i��|D�y�����k���W�mXq�mlq��9\Ě]��	.����-1�N�Y3��6:�w��2���}�{�w�^,��S���
RgƦ����`�@�H2�{����=�?��8X���� X�ȑ�2ֲ����~��@[�"ќ�Y���N�ۜl?�'�l3bh�C��"QJ������+��� 
p5��On6���@�!�"���;�Tş���j�a����S[h�!t!�{G"�f�M��z��yd�iۂ�N4����v
�_I�[Z�j�ˈ����/�����ʪ���?���J���.�x�m�N�k!p�K!p�*�Y��U�:�V�1N=�P�'\��+c�|um��3
m+
`����|���(f��W�������cj��MB��n�촌f}+�)�nb`�9BO���w����JM�*�|+�������^!0a��Ͻ�z�2ô��S�F�uEs�Jg����$�̬�ݤ���G�
8%yu��nGƺ)�\���������,�䄲�Vh�a��m�y�h�[f(�݂_��R��p�0��sh�Aq��$o3t���j<^%���U7Q��D�q����==�!S">( ��%��wd�?����	�Q�&,��7���^S����\�N&M�$�X�=��X7P.�и�s�y��Z�v��'PU�_�S��6��,�G��+ae���{��H��U���h�� &���g��m�M^ߡ���-��씚�Z�Q0%/�J�t\`3�ї�}f�q����&Z���+ЧMu&X�N�5�&^�恗S�c)�"y��%5��;�F��i"W�׋*�g��qQѺX�5�Rܢ��@#�6��D	5�F7|��H=a��E��� &?�+m;v�ܧ_|�u��#��K��b�y���CڽW����n�Cz����n}6�}y���X'/�e��ѱ8,"�FL��i����PZ�O�Q. ߲�M�y+�p�Қ]�w��T0�@���/�Q5ܔ�U"�m0���%�1��3����l6?J��)���l����\̫2�MQ@ͼ)�7�84���mo��R��� ��ݲ2���:��,��ʩ?1�?ΤaV���a��6ʽ	��x!���)[̱�wl�X?�g�b_U�!}|�]h�DJ��XHV���l.�*s�&ʼ��ne-+s,t������ '��R	P0���Ec�x͏}�V ϕHPG,:��k0�?c/�VXF���o���
��c�6Y����l9γ�� ���n�x��5��O`���3HO����S���<ҵ�	b�ﯵ|U��Q5>'>��`�^���n&����ṽ�hCW@Q~�'v���N"�8ك}��v�;q�{{	��?�7޿_����3��������J\ԑ��^��q^�Ȫ,����,�N'~�$���a�U��`���}��Xl�ġq�a?��l&��.ժ������z;�s�f�T+���;J��a]A�\�M6��a���������w��)	A�YI���k�R�ml�C[_���-]K�/��\	�\�L�3j00$���#���O�2����qN=���d_���BvW�N�c)�O���ǰ�|�}�X`��� E�C�C#4���y��c�Gk.Ռ�_����<�t���Bލ���f�5Ts��c�Je�@� �]�v�z*`g/�5c	�Ju�_~�G<5�A%Ύc
�&ua1�:d�Zx�u�g���E�>?���L��"T��+�R�T�g����2Y�b!z�U�m�$	6�}���'zB�MV�_��W�;�� �B����a�|�Ŭ�,��َvv��/։�f���1/����<�"_�6Օ���T����r.�^�-e���:9��C�o'jA}:^W��xe�X�T R��![�D�o'R}�Ƨ9U���g�_:�°{jm](!m��o��r�C��.�o���5�� i��zR��<�^C.␔��������	B���w�,�y������ )��ËP"_?����
�Ki(v������ю�q�r�;�B��	��z�A�Y���{8�?7��N��21	?zd
�3��[�.��� �֫?9t�`>~�;�<����I������S����Қf�ݳ���g�D8Nj�Y�1*Lc������d��v5�k9Y�	7�ɭ�h3'�x�UPMC��H�\ǣ4��az6�����Q�A
eg�4jFp��B�����\��@�=�J�ζ�t���ܽ��������3`��]��ϥ�t����4*�'�aBg��9|���_�@{���(=2�6e~�U� J_(+iK��~Ag|IP=y.�?+���s���`c�-I+(U�'��ȸ��R
�w+�ʂWQ�PB����c#�i{� �S~�J�'���qu����"�� �q��36����85��ǆX'��Y���7���K��:r5������P��&����0�H���J�|�g�>�c�>Q��|�A�9�8��NP��9�Y���¹��O�Y3���p%�u#bZ���"�v#�%�/�0ljs�̌�x�Om�cF�Յ�fN �*61����r�ݗ)��=�?"�6��j���N-��s�[�ͳ���C��|�.�~&A�L)NqN��wq�t��4����oC+�\��cy
�O�>�_hw�)�������})�4����TO�t.�W�.���sS��g��XGƞ.���H��p�u<�ڤ$���Ő�Y�g5%)�-�'N>4V��x�F����ܝ��}�'̄M#�L����-��K�%�|.��Gh:���-s/�u"���0����lNjV�' -����@�bH�K����݊@'(V�$��i_<\b��X���S*�*�?�U�[�N�� �z@�{\*���7�/9�ǘu�&����{����!��x&D�kː�
"rO�^��]w��5�@�ԎA�j,plL ���2}��t��>���5ɞ��i�&9��o������"�^

�⸦��ȮQ8M��%�k�m����mt�&NhM��ef�_Df�z�(j#
����	*	��9�|�D��m��ҧK��б� ��.m�L�쒏���BE�o�29ŪG�7H�fU���k�"��9i�*y�KZ]Ai���x����gl�m?��5�O�����#^#Ə�G��w�����F�YM�b�O5�F�0��E��E�ϧ�D���h�j9��X���硯�ș]6L�I�|)���@f��Z�AW�|�����	;kM����m*��4��ó�z9��e4ʹ��C�!�շ�ruIa|&��@�`���nT}����jB|���r�������~OH陭��$���a�:���˱�׌�-C�F��[P�Hw-�Ԇ"JI�2aF�`�	���.X	�x�M�rN��Z���"�ls��d�@bU�Ƀk�4i=�~X�Y�h�G�Y�]�k
Ѽ�cf���7$ }�9�4���+ض�Q��2�<*�E|W0��b�6���;.�*v<�EStV�Y[�;ע��.b<�<�ܫ�"��E���կ���FV�| ?�RƫRb���斕��hAhi�������G�xK�ZX���B \E��څD�+BDj�lAP����&p�'�Ȝx�Ө,a�):�q���hU���T2G�%e�N�Z���F��?�s�B4TS�{ٕ�V�G�*�e�ltx��	4bHxe]��Y�7xy���Id�R��j�Y離����~��ǅ�*����[��F��=	i@zA,>��w�&��N�4�����[C,���WH�+W��Et��F��ἑV'��%�+��c����%�C����(�玄���%*��gn;]�v��7qPC
2S��6$�|��d�QN�;7�-^�T᝜1���\��?�ٴ��e�9�D����~n^�YQ�3���;�~�����6`Q����-�Sղ���">�H�.�i.uz�
��X�p}gT�^v�貰y�������H�֔�d7�����=ˆr+?Z�uG�����j�}pޞݣ)��8��gXK��^I��/�<��Q�/���Zjj��e�|nX�'�V�D����Ñ�M<�3=�{��X%|]�l=��W�,����^z��4!�������)T��ۋ�D~t{8#GT�?�WBs7���ʘ�a�D�z�u�d�H.������5��6�Df���Z��͚�M�� +5�p!P�f''��#y�\`�S�!�>5����;M���#��a1f[�����G�_��Ȗ�W�<r�`�!�1��
e�:�G����$����Ƈ���\���!��C�^W�#�Xhck�6ɾ���R�}G7竕�ֶ��2t!n�_�*d����]GF�v�%Y$��-�vr(}k�%����IT'X�ot�͓�q�t�K�-����S�K.*��p;����?�ϵ� ��]v��k�cĐ\�������4�yRn�}�=Q$�uB��M��������xH�U�5�\-d�GL�l�	��g*ԗ`��!(27������kjܚ�¦" ,���ߗ�f���z ���r5�p����i����z6�FW��< bOGf�hP2�sP��Ā^5�dn	��{�u�o ��Y��	���@E�"@��QB"�ζk���CG��i��˕`�ګ��_�j�����֟���AO>ATˮgDb��Q!ߍ)��'H�9��Q �r��daaE$���)f5��Bwi-*%wI/I\��+�D�-�����.l.;�4�y��r��L�4� �F+�n�	�vy4/��m�S1c����ӏ��&��̞�U���B���~x���������V���Kݞ��%�Ľ��@�or��ed�W����B�w�o9�:��K�:�_����qՄ�G��z�2�V�+vxEv�Q!�����r�ێ�b�9V��.�La�(����cz0Ta���G~�����ݟ�/o��}�{�<rhw�|E..x����5����%7�V�L�>{���:2��Y��͆�;�
���̟��QW+�[��`���k����N�S��~��e�I�[#镃�bz��q��N6��x扠�����J}�Fn	�D�G�gQ"[z��p���)EC*e��Ƣ�2�˷��%'Q�C���K`S�%a������Q�x�<�E����uקw,k��'�Yu��nMh�m|���p�;42~�7���M�|�̉��4�<Y��s�����xŌ�Q�Q4�l�:�`�8gJ�m�)���������^�xÓOs����Gq� 6Q3�{���׭�}�� d�8�f�$�4$�t�,�
��y�
4~��|�l��[q�����0\��W;>�ՆY�5me�`pg�~����q�o��~��6����z�lѭ��H�I��I�xR�����rA�KV�1�߭�{_I���Z��а.���H�N�Y�����/�����	Q��GƋ�WsLH���V�93�L�o��8�AKZ�U�P���C�)���ɔ�G���F�C��\�/�+������s���+5�p�̐�&�鲞�w��m|��@O�����)��z�g%E��U�'�쁥�l..�t1�PձF��B�w��@_�1�UR(_�g�yej��~��#`;�*��=4͌��P+#�Q�tp�6�ciZ�7=�$��!�CR��RX;-VE�N���JU���6T�
��V�����_	D�\����=��ZQ[����'�T>+
�N��nkc�
�pd���:�fCG����8��˩�T���4��Xy�ܻ�2b��M��G�8��J��\�9�{�{�4{�&~u��uRk��,�a
QЖ����jQ�Yf�;YvK�-�Ӯpt��y�V��/Z}�Ăٞ{����K�bu�x�v3�AV�kY߅>����)�' "C�s�Ć$E��'����*H�rNnZ���%yl�P޴X���J��h1B5-oS�t��f��C����z8�
z��ȡ���8��/'[邃Bta�
~k1�����=ޚ�,��C��� o%ʻ3w�Ka;��7<�f���l�ԝ�|_���#�sʶ廹�5&Bz1QQ)��zWeҷ<����ǃ�}�=�;�GS~�<[��g�t�g���ʹ"����'�]*�C�8�hi&�X �/?R]���ݜ�I�e<��a��<X�}Fh�>m;��6���!1�Ji��s��ll�\����X �EH�M������YE[@��Eɘ61:�b�1�i0@�� �*�)`BV|�@�� ��Cn�%-@�H�̓祡DbnQ�<��r }�04�ak����t{R� ��+dV��!M��2�u�"���.�Y05�Ÿ��q�'}h�,�Ȍ�tΈ��D�B?0'}��-�
�6+Zh�>X$�6�0;�n���5�b	���޺*�����5�}>��>
k�=�$�Ċ�^礒h�ƹ�:�j�pU���ɿ�q��<S��UǁQ\{��SDY|ϛE3Ea�3E���]Ӻ��h���GĈ$9���Y	��
��jyo?S�4sI0��k�w'k�g�Z$�_{�53=D�u:j��VC ��e���<�_�k_�vq�����Q�K�^���XQ8lI'	I7������ ����D�&u�w�%�.-)�� �����Gy1���*��w�>�2�T��{G�Ωmbx#��������1�$i�*���1vy��i�	WG%<�f���J�b�WˢV��S�.��?��M����:�d�Д�t�AW�	[�e2���F�e����%�3L3����$��0 ��>%��S={��ʥ����:�=��v�C,���E�_�)��䭭�p���ju�EA�١�����4�Qt^]ŗ�d���=E��u�5��C��}UQ>.yb|E��f�|����:������j��\����=u>z���,~>/����|n�I2�5��t�����.�UJ5v�gEeG��!�d!d������y��&Y�rK�NP0��C6R��L��=����A �9�VԌXTyU�
�ɼ�c���?��Ҕ"�nO#����uMx�K�� v6+�z��rZ����T��9}j����C�oL��bqA[�Vk�u�9���OA&}mk��g��Y�9�E>?gk�͙�����|dTc������S\���.q
I��c-lc�4���}q>獦���>S��mpz]�A^�@!�H�
�\ս�33�w��4�i����"�y��d�eP����0^��J�2#wT��u��rׯ����#�=ux k����<fg�MGl8ⱱ��z����Ү\�OJ��R�cS(���C\�`��9r�sщ��)�h8x��@B��*eZ4��v� }�$�)�g�����}�DHB#�PQ����oC��#j+��$�uޮ���}]Ӕ@������ٔ��e~��(�O�=ɱv��V��x �C�3c8L�/�\���_��15������~��G'�����C����w����nr���1f@�>.�P ""Ŗ����$	�����F���^5�:	,8l�͇��uD�3��?���yO��W1�y��!Y%�اR�@��`���8=�?�z9�����h���)��1�'�Q&0�� �\֫�쉤��c�TK`hO3�ݑ�jk�/�d��7hH��<
�Y��C�'�|��0��l
�5�� ���S�#S+Y�Z;̻=��Eo��]hBɏd1� ���e�;wZ�VxX����W���>��O�zW{�F��;�g�z��{d��Խ����9z�Tst	~�S��S-�nb�ҁ�������(�L�J_}���K/a�Z�n�����9}����)�E^Y�)O�̅�������Hg�g7{�Q%���b�1�A}`o3_@��V��Y}lG������|YV*"�l��]�U�
�L�*���+xl�ާ�Q!��Z�F��L.��S�AK�Qv'|��UN�\ac' or�p��V��Um�DO���C��!�G!�����ǂ\>r�v�,TT~:�k�����Vw���K��r��χ�	*!�I�I���<�b�N�5I�g��g�"��eo�7l���d����������Sv�}��tq�8j�֦5W�LN�!p0hi��s۠M���9��'v�:%��ٌI*ĺ�. �)�(E�m�X`�LD��kK�E�F��V�
W��_��W�gi�8�C}� ���Z��	���L)�B?��&6d����x*� B�p�>S������5bs�"�8�t6G yT>A�=8A$�����n"�Z�!�%O��s6�F",�ː�}`�"�� ��e����\�=�ܭg��2%{%~\�J��o+"9Uܾ�� eF�hR�k�DٻP��i-�~�/J`T:ej�oMlwI��qZg���d�~�Xv��F \�<J�%ȇ�Ƭ4X>�b���Oq�,H<��3�(�N)��R	��&�h�)��zQ:�ON�����x<.Q�0C����og�!�	G�"��꿫X��g�$"s�转TS5�!`�f�Uu����Bi��/�۸=f(?c��^�f�tj?@¤Է�Ls��(\0�[�#~�/je�2��!�R�l��oE�Nv>����(����i5�d/L�*��֩�L�F�:�5J5�@����$Lu��!ٍP{�ݽ��F?c]��ͷ��1ɧ_rr{�4�R�U=I��<�5�QN�`�ۡ�϶���h�C���)��	�~*߉)H O1<�!8������������C�ꏴY{�Xi��D7���T�ER�n�"_�Q5K�I��"�?�Ng>Q]��4&'j��B���Y:V�f�v@�_c�0�A �e�hd��:ؕ[�]�'���|�r'1N�SCZ}��'��FT�Y�&n�oV���1/f5�=�<��{p��Z��
�TmgD���1�]�F%���00�~%�����M>mG0a��@�������w?����q�8��p�֊�ߴA����@�|�i=j�`j�q�I��t}1����v	�-Y9������i��2���c�H��MaIQ���޷�*7���u6n�,�}��h���<���~�b��z�����Ap��+��4�Vh��*�ޞGzaX�ɟ�M��Yzt  W/F�5�Dj�eIKG�����a�W�g�p�'�p�����e��]��/���g��qG�7��&��T��%Y��r���2aI<�Ol@�c#PnS-L��s��ךRs��1#Gb�Đ���^8����Y�)��q��<�!��7G�*�/k،�%y����|o�9�mz�5,C`� 4��s����4/pܼ �o�}��t�8\چ�����p�]���((�89�b�&�x�{��������S�W�x�:_�H��EH�p"_�������v+����w�8�?DH� %��h��w�FQ���[E��NJ��Sް�D�#�Q&�|9�%EQ���.f�2g��&-���y�2�7���Tj`D.v�\q���p) �,�l��R��}�C��)wJ�ۣϞ������K͔��W`�d^���:
��3�Y|�_���
�CN�ZѺ%�zA�<�{�8͗]��3jǺ(ZΝ-�E0
���^2���.�t��I����&X~��
xt��8U�1���vU���)%��r����R�FiN�b�K�zR~�# ɅRy����lt8ߝ�R�~AB�~�v{O�'��L�2wH�B��|�@�T"�[h��`���fA-E(����*� [��#�󉖠a@4��4I�"Bm�@�\X�䄄~Db�bKb�����N�	r�$��À���[ڢ��U��Q��#���u4硯��d���(Ë����{+=�wQ'���Q���|y�@n�����W2MO�Xԃ���ѽ�M���D��ͤY��$L�p�۔��k �^a�®�$��?�pKsK��z���eʣ�TrB���v�z��)^��׋p��B�Y��.����������	kx%N
p�� Dh�i��D�<0���l�&'{��@ݥ�Q�N�c��I`-/� �?x�b��<�:U�>w
r��
��`G,��4�����"��,;İnr��R�h/u �u"3Aǫ�@��T^� �k͍���d�NA3U?W��o/}�LS����i�����uF��:Z�nomuK`�#�y~P�#��59ttd�uv�g+a�2��9�6�-�ٞaH��������.i6@˱�Q�F����܁�+|2���יp�8��3"t]����頛3GP��#p4�>��gәF;mx��X�|s�s�G��@K�#5�Oz�"�	��lXد��.�G�Kk��-�����`՗�V9^h�>"��$^u�_�4v��N�J�YB�<Eu��������˃|�֮h豗�ī&�˫3ê\�exްrtYDh�����c�G�
&7���V��6u���k��Eи~��h�%�]�!�K(�����/Q�[3��� �[]�EI���e�AN�ք�Wa_Q;	ܠ����W*�vK���fO�.aH�����u;{뉒X�
�q��x�0d�Zu�T�'�����Y:�06���jn� �$CN�
�-������M>Ʒ��C��*�Jچ��������$ҟ%(y'l�C�^`�5[����t���Q��\D�\e�/���6���xjP��̦�V�)�/�R��ᤥ��-T���C��p�$Q�Vp�q}��DI�D;.ej�|
'n�ǎ��w�>�+�GT����J2F���
�ӀnlJ#E�&|�lS��>@1}׳���m�㔶4�q�K;0��@vФ�
3ע~�D��ðW�_���7������ɑЮ�i��>e�^Z��b�ᘗ��2U4�ɵTe<9�wO����L�@�S}��e�)�����GZW3��AB���
�Wz�jaȂ]J^�
ȃ�߿2{�����Ա2�ۏb7S��"�}�k����E���t۫��"�U����.��$�9���f�����Q�~��@,'��˒�ɢf���ݓ��$Bo��>36;�k�����o��s����ޓ��5wp��tp�`s��b7ˮf�P������xA�n�fC����8�N�3���$as�˱U�9jP�Xy�7�@4O0����hB&`,k ��q6uq/\]���9�g�6���mM�4
��(��fL��.��
<L,�)�~�i7�呏h���v	n�҇r&��[0_W�l��>��CA�@r��6��m�����:
bX�3E�D]�ҁ�R���ҧ	�]�U��,zø��*����$Pi�������{���9��<@U�c�*�')��(K$,�q�nC��W�����;N.3��gg�(�.�`��b���\��m�
̵�����2d����S"��3�
�U�+����:�14����nԄ��6:���!A��A����1_�*.5�&�mR��?Fۺ���_���]=)���$�9|M�{i2�1z�����҉W$q�a��\�����l��c6~����fSd�^������9MU8���	�lj{H��������l�Y J_�x�0 ���et��L�~��1��3����t"���Jֆ�Zjeqj#�L[�"�L������d_���G�[��&�&D�yZ�}O�7���{s�����͌,l�j;b��ԍ,���O���ZT�Ac���c��R��t�*D=���7��W}I�Je�
+��Ʋ�a�&�����{�y���� ���S�R�-C���w���2Q��A��^u>~�:�L��?q?S������-�QZ����
N�Ez_R#%ScKr}=?�^J7��˫�q�M�0���s���D�>��ےT):�b)s���#����	t����V62p�r��r�����3�
|�L2_K2Y[F��$��p7����������<���bJc�4�r45ͣ��|�a��|R �p�����l�<g��i��ʉ�x�ԕ�.;.�
l��YFwĂ ���D{����
�g�O/��P�G��=�����o���0� �b�AZ�!�zR��'�o ��E��oi�Tl�o?���
=�B)`�I�ɦ��~9Ņ��>�fY���I��k$1d�M\��*���6n�9tE�H�lEy�X�~�=��T���µ�@;'�W�S��AF �m�2O��5)��{����� �%�3|�3�ց�=!CI.�W�����qY�k���ߤ��wrFP6q���]v������r����y�^�MHŃ��zjI�$!V����$Μ6�A�4v�CT���
<�e�F�h�]��]Ip�B�Ց�ymOBi��I�78|YsY��f ����Ԣ��� ؾ���&�e]��7�|�I���%�I�α��6�F0s:�n?r۴[��r�=9A%Rm�ou8��v1����+���R>���� ���c�������G�.��ߟ�y-zbMΕ4D!ҫ.H��x��˸5y.�	+��Ң�7����Aj��4\i!]g7,7��_*3���x�sFq`�&R��%���#���[��c?��]_�",�I�ľ�k�;��I�%-��Ȕ�q%���L����o��t #��e���R.@>/FL���qH�$����1At�9�(HS��{{;��Ki�u<3������(�:�� ��X��i�Q�|R$_g��)_�D���-QZ$�.^p�fo3l��n�� ��Q��7��K� ,�[�4:Hr�18���-
ܬ�r�~�E�?t�'̎a�R�uL�I8�K.�"BFF�`��. �����s]X`�0
5#ɣ�T���c��_<�B���	7d�l�eE��Z��3����>į�oô_O�4n�͆��d��<dh-������m�6��\(�������)����a��g��P7{ex��*w��!�0������lW�0eO�p]��^w��+)T�y�J�_����>4������l�;=�gR-QI�{�{��H�[�?e�:w%ĥ)����K��k(gȷ���x��"Ra��6á)0�w�H��|h�W?J���+�lu�0��m"}�=� �j�W=��}a�z�ܘ�����p��gM�����b�?Hῌu<��t*h��3^ʠ2uB%}ux"�Z!}�J��M&�E�@bs)�v|6�v$����� ƈ��4���{�� s͡d Bl��� �$s7�B���o6꣑��� �@g�����z^�Y�z���N������}�<��G��F�Eq��0cm�z��qJVy̢5)��Nr��7�`�˾����	=�ס �q��(��g�zi޺�	��RI�s�)�5�k�reCc9O��:&݋�q��u$���s%��^��������MF%Oir�> \��p�����ǋ	d�z�C��*@M�ڕ$0b�4S�oo���*��wV��w�*�O�}S�<u���ؗ�,�#E�t�i"�o�Zf�N��5�-&~������&���Wu��8�5A$gc�B�g?"Xhd|�\�L��O��Vo���.&�@G�J[fB4�A�c�8�R��I-PHq�₻S�w�Uڕ���D�k���ձy�nt��j��I���o] ��m�zY�ʩ�I\�g��H���O�
#qV��{�qKWi��lLg
 s)H���Ddo�~��ey��Hcf�Fy`���k��~j�� )�D�ʡ���!ĵ�#����
�.��~��)�4y�ȍ�l_0���*�o�H��=��D�l;�ٷ`gK��tL׮Ҙ`~-���DoA�|N7*M��d�l��K9�Lc��Igw�T�JY��<��Q�)Q���4�d�?n����w�x2yx��bS����i�:FY���1�����~i�T'�)没���m9Q����<���-o�pn�����>�$�(l���X��Y�E${[���[�#=@4/㷇%4;��<|�%�8�����&ra�(�+y��[U�!�����JX����~�+�t4e�3��p���<�����ow�wCG(�OA�#Ā�S8�L;Z0R�%��oiG���ĻR��畴�`l��D�E���S=l��k��Z̦2�0�!��YU6NL���Sx�T��ͽ�,;e G�������Eq�� >v�o-Z�*2:o��\�yn7w|��k��`�����iQ3�(��B��A�M�К�>-H��H������gd�`wp�T�U�=/nM=��ι�三M����9A{-��XF�����5�,#r�$hZ7됞� �a,�P�z��Eɭ��x�r�a����� �&��E�@M��;< O8f:/�Y�a��mLn����Y_�K�^sx�]]�G�mQ�����#P̜8;5�A���t��$(i���ϨG��'
���	y���5��Q�M��2��J!������u�h\g?�O�������#F�+��V��a]SkKw�D,�i��?p[��|�N8JD���� �1�F���E��3���l�s�� $��0|�(z�UJ� '�y�Y�؇���S�2����gc-��+D���g����$�+���^�E	�B5�D�E��>Y�� �f�S�B_�Oː(1Q��[`5�ꨟ�}�P�}����~��M��t��i%�"y!k��*iÒ�gX��z��'qp5��q�}�h�Yc><�)_����΁�>X�_F@i"AH71��/��F4��o��p&���T����4ZẰ�E�"�5��T hRe"��T�QX:]^�Xe0�3���[�Ԯ�h���e�ws�
(�)G]��Ӊ�mOWC]����c]���E'6��\��|�m��j-��c��w��2��W���:�*���(��)�a�����0~'�?���=�E$P� �sd��(/
�����1���eZچ^ ޚ��#���>׌F�
��!��ȃ�M���H�3M	���rbv��vq�B����5?�V����N�Ep�)��A�{�4ő�V�0M��H%�&,���J���1<�9I�g��kb�5��L+�;�6�[5������&�bS����6һ��I\�1��� ���ir%��B|��M�n�*�bx˩�n�_ȴ�'U@���!B��LJ�\�(���I�X�j�c�^�+��qc8���o>j��w���K�84խќL�E���j�{��7��Ȥ��,'7�?�4A��7)�Nt��A\0�2C��BWgD�lF-����m��(=���u���ɨ��]z-�6�/z��e��FK��"FG�pB�*��E�f�����B`�
����I�p#�U�	�FUHK]o�Y�P�c2�s��"z���D�7|O�ť,Gu[�@�����%k�ε)Nf��4)�G�������yo��-�@�G���֐����O_�C�}���ƦXԐ���z�˸@�����nUy�A~��0&/�X!�:���-��J"�qA�I'c�_��9?���>�"�־�+Ɇ�5c8v�յIP�F^7 B����:��o��T�1A�Oh���(6�Ŵ��B�f[������s��|,������j��J��P�gD؜���B�y�"���aV�հw�d�>��_f)tc�H(�Lg��מ��?V��x�_�B���~r��S|��C���ŭ�\���
7�n�4��
ʏx�P��-�g��2��K5!X�k��N(V�D����Յ�|?W!���T�a��:1`�����6��Ce��	��S|���_P����b�.}9�6{�-�FI'�W��@Mk�,'�K���/(H�s�	���,xQuZ������I,3��$SF�R��i����bA�QU�	n��)�xy�½r�g6��o�5�w�s�2��~��k�f��X�P�\�Y����,|�hv$�s���A?���OTL��x���O"�"ރ������6�TԊ3M�v�v#��մ})��=�Gc�O�� �؇w��E7L#/�v�
b�%����PcC���9�T��o����Ka!�����u�z�Q"g�A�g����~&��Q@L��e���O���൮F��nhi�ޅ�����mR���j�� A�vN�3�U3|px�)�і�[d[p�9oN�7V#e`2޺h],�K�)� ����ggYӎ�a�p�@�Q�� B���- ���q��cq(�Q����]yڕ�l��=iʸK$������i�r��	<����
]�#1�K\)���v�
�$ffy4p~)�O�I����t��Cϒ�	�
���},:8�wGnY�P�v�zP ^+0�X�#�汀��2aؼ}br�	��S��yW}�&�~�;!u�6@�H<j�h4g�������RA��כ=�ZŨ�� n��H	��Q�e���4i�\�Y®��ۛT�@TG�����Rs�J�D�x�Vk�$x'�����Ϳ���۠`����J��z��� ����9��j�;���$Mv懅�~���̩�&,`*B��L�����|^3ST8k����P1�w�(XJ9���*��UW��:.6Qk8��<a�_L`ػ�#�0g�;I3�j�2`ؓ��s�� ����/>$�]�帑K�Y��g��l�^ѯ�n�d ��B\]�h�ո�~S�&�_u�b�����4����T�bw)5���'��ϫe��<���E����j��o����H��.E80�E�y��I��s�D/Ź��	����p+�AJ/__� �q�%��}]���Ъ������6���T�~5��3HҖ�o����s�[���r�	�����U���@vM��p$�~�O|Z0��9Y@�� �ϊ�7/��t���v@���ю9�P���2Hc{PY��9�*�L��l���w����цr/e(�Y�dR�f^Wx]'��!�޺0|�+�+�h�J~��q*P���s_[���>I��1PW�4�\�H����
ؒH�Tw���5-q>�4�'W��6ik����t������@]%�QV��䦘�)º��I�Q�|�'���́���zL���D��j>�����e�����h{�P��S�/���R3+r�%�Q�$��	�̊�l�#Z�[��U<��f��h���!�Ս4qgm��Y����<�ј&�TK]@���|[���Iy�����y�v9D��B|��5�4�X�`��&���o�J|�[��T[��ƋAv����K���z{B�C�E��K�8J+�z10����oT�b˨��<<>���;�'���49a6��Y`u��W�B����e��G�)��!�CC��5P0�������������z��f�O�^K��,���G���a����Y����ͧ-,�	��%��!�w�v���2aq/<�R��/s~����%�d������C���'�� ��������SIdA���՛�(������C|��JVxٷ_��L1V��:�}�����R�����ղi0��g?j�0vI�jΈ�I�`H�ae?����6�̔���(�h��vxЃ"Q�{��Y+3��9�`ϗ��*`w�@�3��'��c9���f%D���U��-R��F���Q�B��m�^�>a�+��-b�@�Q$��z48��B�g�%���l��,���IAz}��v]�)�S�G�e���h�cA�&o)`�)���C@ߺ��|�8Wf�)��m�k7V]�o�z,��.Ά���`m��Z�E��X�Q�:�a��{1|�������砰��H�*8fZ*֢�F��bk5�Wɶ���,�{�bk�}�w��0=���e)��E#���|QF9�&:���|��U��F��U
��O.�f���eR-)������;3���%� �O���Bv=X��x��^�C��圠,�A�j<S&$�B��%)Ng5��Ms�<������q���������a�
@P`��]�p�uK]Ԯ�����+�6t�������Ӑ:��v̓}ڕS��D��j6=�= ��}AkJ���v�TΛ:��kS����HmS@���!�B��e,z�f}�e�;�h5��`p����������g�*#�����9t* E- c�����K�]�M[r��g>�ڬ�Q.]��V�11��¦T^�I6k���$'��Uw%�[6�Z; �'E�B�����$��l�a=�U�#���K��af#".�<G-[zG��z�:�����A�a�u�ٗZ>�"�Y�1�oM�]0˘�Y@�{�mJ��u��dS\z��� �e峌�t��D	q�#v��,����aW[��mx�Ln�L�+@���f�r�l��K�b7�R��1�+7���,v߄nQCKڜ������l����u2�U���@n����M~+����z�����<Ѫc�R<[a�-�Ge0�U��>��I ������	���c7%
�3~�Vx�l�+!�R�3�@bN��E6�J�_Bo�Ɩ˭�m���3�;�*�1�j��܁>ky��%D:��5�3�alUe�!w��Q,�ÃؓK��U�r�<\�Cg�s`{�mD;T�N4�x�k�F����o�R-}1��"-'��H�o��8��8-��]��v�|X�w�����a�"�l̰r�5�������������N2a�\�L� s����E�?�Dk?[������PFa$��ːUˊ���by�?�� P��O�x�Z���9!ⶇdp�"�f���aB�����<F�޶ �v�%���T�������2�5��S��?�����7<��3�U$퐇�l�� H+�����}�y-3�	E�IPj�!�����	/uN0�DqP����p̂��|�����MS��4�j>�9a�т�n���;��v���4,Wq��=\Wb��Q͵6��v�F�;9%�7|��P��&��I�-��.�?��\�*P|}�)�x1u���"L�2��MCM�,�������L�!��oOދS���vhG�j1X{�Sn��}I/�0ۗ�.$�i��@ߙ�W�w���K6^�e73 /A8��?�tJq��1�+�����gg����4�؏}���f#s��`�Z��{�k+�E�tJ������`iJ�`񒆙ZD3�\���^9Y�	��?TE=}<��	c޸�w;��w��W��&���+)��wU���\e�|�!$���3��[��M��մ*n�]�����rW%y��8���Z��6v�i5�	o�$�����튄g�u��wI�J�0٢`�&��5SU�a�5թ�#K�2��;?8��@S��ůkB��$Z�'���&FHhs:N��O �Gϝ_
Lk�|�Va|�#'�T5��c��4G}�&#Sۃ@@�R�������`��v7W�T�M#��q��̀�z�ߚ\c����J�~D(�C�4�S��NN����*��9�b6�ů"]f�P��f"��<��z�`��t����>�%��`hG%�` �$psE= vE����L�,t������|�Q�A�WM�q.`���Su�F2��zG�:���˜I��i�@&�m���(5�e���]z�.�n	�=?\=P����&�2��R��ԛ� 34�-���YL\79�𪟨���K�	�F�=���B(�ڂO(�6 &j8�j>Á9ږV����f�1!I�dy�E#�#������E��Z+��z	��"�������ٲo#L��`rDG7�@�a�Ŀ��2D;#�=W���Y�<�o���m����$fF?��2zz�7�1��%q���1x�&Dؒ���=�q�:x��G{������}M��� �E����T��"��^~�%�3A�8_	IpGr�~0	�����V�z7�)�!{���m�U~Ǿ��JƭW�7��n5�̃BQ��ǜq��ޱ���e��d`����
�'�/�����?Q4��i�ML?�+nf�IW[��EDv�aj�+�ΈR�Rsm��2�#�1����n�E�AS%�x�~�����|ￇ�M����ޜ��S�|~����=���9����]����b�%��d��z�]fB%ĸ��|�5�C���뾧J�'�*��mU��Hb>X����<����c�8����^@v��O��Lo��"RZ������G� �rPh���V���nC	@���:�������'�62��]���k����E�.�R����Kxk*�$��)�H1�`$-|3���^f���]fd������ ��vߗ��H� ��qTΦ�JC!��;����bV*ĕ���,�ܖ�SԾ�YЙ.��k�:LG+����9�G����h@3��Bj4U���~��C�N�F�w'ئ<��9T���Dc�t��/����x�����<,`��|��~�[3zg	Ad#%gx��=����xE����~�r0�������k�'B( ���=�\��6���f�<F�Db�p�a��\O�㜁aA�1��栃y	]^��I{�
8x4
�cnͽ����͵���f��7�������Ą�3ˠ�FΏ_<�$hnsҞ��ʦ��C�P��@\�@M���T��ـ)_���2���� x����	GO���w)�%��Yn� n%$R_�8��;<)v(�}>ᓅ�ﶘ��1B��dc�i�C��o�Ú�P��?� ���F��Q�\"�3�]��Y:9�<�:!Ol�i�[(k��䣠_�Lc��9��Mu k]�t�|��(� ,�~9�~���YoFm�-��ý�)�$7�]p"��0���"���R��԰a�=�N^ j�,҅�F�M�\N)j�~�M��z��������'j�����O��_�yL�	�����h�zd���j��Z��$��������?M��õ	UJA�A���m��t �c�����V�Ct�"Ẹ�˂�..w�^^�7�")��T���d���%ǋ�E�w��&8w��S/���R���W_�+��p�w�t_�8�̌#3I�WN�F�
�\%Py�v-��~��]�w�ss�8a\�������e����ݳ��;�c����3s����"�~.����g��*���>e��+�{�����N!�]>h��фq`+��pE������{ym��ο�@��zM�n�uu"׿O:S�[WpSV��Ui�*�_�Q6+��#�ޣ�X��TI�(٘��di�/x0&cH�\�{�R�,����֭ڶ�� �c�	έ1 R��m$i�ߍ/���}8G�z�v�?vHíA匔���H�u�I�mLw�iybs3�<[����;ZN����¦��,h��ABAK9,��x����#�]��?��,.aq>$ɇ��:M��?X"��$��V̩�a=�_�܃��i ���t�(����v=_���:�i>��^'��z\���;?"�j
:����'�#�51�[:�j8o�>�ݡ˺@�9��S3̧J��`���i3��G�p�!�	(�W����+:}o7cG�qvPy/���S'�-���/�I���&�V�ڥ�C��6�֥^�����^o.���X�F�|`T���O_+'%��X�D3��]x�|�c����pΊv�I�� J�*�U��@C���@�@������(�
�+����L7d�4�K��]�]�ь�!����/��k�:�M�޸U/,�x_<t
���!���Ͳ&V���	X�q�OV� �=p�S��g?��)��mՖ��LoP�u��݈���5% �غ�1���0���7�EC7VG C=��?�Zݻ��Z>�>�ILv�Ye�m��h�HQ��?�@|�;�A%�0	:'�a�fǘ箉���[9 �i�Q�jc�iR9BT��M1��X�+^��ν\CZ������2CP6�j�D���T �{;)����G�ۣ�Ƹ}(�V]��\����n�Bܩ�.�*/�IN�uIka�F�<̕x���S��ܐMCϪ�x�r�R��s6��3(��-�2';�EF�A	����l�0+f�v���2�[���<N�\�����%��*�A�!<��"�����A�*�S'�D3g�h;Rb��ڥ�����.��1o� �j���^�7\kK�Nw��WC�1�DmYslt����`̖>	a<X�ǓE�Qd����Ų�C(h����JB��'��P�������g�
7�-�rly��}�^�􏁍Fu�vʬ,@�Uv�@jRRy0��.��zrSs��hG�.QͲ.Lno��K��V�P��U����{�i�ںD}���Y���SW,�c��$ȣ{��L̕A=�}�3\-J�ċ6;�[���ѫ)�hv�G�.������gڇΩk�01I�E9�<��
�߭ħ�sYK��z�����*��ȑBcl\�M�CA�C�.��h�{ZxbȆbFbQ��V���)w�7�}jL%�3Dè�U����#�� ���;+�)d���G��	v���mdS��߃���J[�	���AE�N^)�`V2�� ��ü��w^[����![��+>/���D���7<!(���H��<�9jG�/׵%ˇ��i=T�> G���T�;Gޅ5&yV� Ú[��)�~�uQb��n8�g���� � ������驘���.�7���-d�k�����F΃0�~���"�������*I_	Fq��ʣ6���8?�]�.�A%�z�kuk1ĶA���)���	l��e��Ҫ5Pp��1�:��	]�c°3䠛O�}��Ѓ�O��	�9=�l�^���D�-p?��[C{�r�V�yv}Ǒ�lc� @�$zm&�)��bU���C`�7����7#z��%�(v{u
fP �'�B$s��������
�*���`a�Jjb=D�y'#:�e�4��3L��D�GG44H'Q[����d�Tg](eMS��USa�'/ �+��S�b����:�)�S7�*�К�Xv�;�^��^�o�Bd(�xVĠ�N�|���z����0+�=��P����'	���E ��i������4�ZbC���m��fL<іhp�zp�:�y9�I�Ӄ�NN��O���~z�6��+��oi39�]̓3?��ұ[��E[���m.��rB�5x���O��e�����-�R���[�f���T(S=!����ӕ�&$�s�C$iQ//Ġ[y���U�ez����d�֞S,-8�l���ハ%U��91�/^T p��.wP6>+m��]hP�v���u�+�B}�(��Q9A��2З������+I����%]�-MJ;r�l}�������=����hm�:8̹�*`
��|H�\g+}�9��s�I~ׁN_Z׵�Ry�\��k��s|�H�B!��?C��#�z��=g�ܷ�v����n˰����F�ƻo��Ȍ<��2� �Z�&t2+�����vl��m�T����Ů��;
�lh��U����+D=��}��aie�,�R�0������gn"�8���	�H䚲��x�6bZ�%�����-�,]�wn���&��	�ɠ�>�5"zŧ�D9<]�߀��/u�D��'�2]��n���Pf��̦��q?��,��Z�$��"4���ފP2�>�q���7�����%�v�0��<,��iչ��:�y�7�I/�
h��F0PO]TL��yĈ�R�����l��v�N/����R��T#:��4�f>nL�� �������r5'��>uR|ʦ�n����_�ey&�-2����-mfv�%������Y:=S��_��w�Gz :g]��\D$u����p�\v9�}.���k�hB��4g�+ W�.����>
���bOU��e�AoPs]� ���ѳ�Fk;��Z�gv��-ÝB����s�녩N{������r�5$\�M�$�W�����6��_[}�/bk��
$;?0�"�%�����XB�����G����&��Zc�ƀ� �[��]�jiӘx�	m[IM��0d�U%��YuS�^UTҒ���L{��k�4A= w��,(��39t:=�l��^������A#�����9n�Le���Nn�G.�Ґ��q�Sl�����k�A��N6,5��K���I&0��/3�Ăp���dst��l�qO�5��w�(t�ޟu3��b�ơ̽�ت;��<�i��i	漝N*�re0g�Gq)#��f��ĩ)w�Ca	e�L&�ʐq����#R���C�>��)O�5�D�@;�,���j&�f\q�c��7i�3 l�'?g$Wݝ�K�_4d���h��m��I5�"��*�ڶz��I�����qA�f�.�Z�XkM�k䴀��r��a�<�(��Rhd5n�޶hJ��1}�J�~~m:(��P��V3S��}�9si=	�9z�hE�'�S�]|�B|,c3LkVj�޾k�*�m.`��I�ź���w�6ȁDQz��t���bH��'�uD��Z]�9m��S��؟=�'zU��qw�-�IT�!!��CV!�h��W
�#�W�N��������B�e�%˷���DD[�j1��*��2\t΂��q|[����B9��?�+�
ζ��.���J|W��M���E�����=�]�c7Q�r���az��(�~�V�]��=h0.Bw�X�,?=F�)�z��S�٪��ĆX���*E��~U~���q�s�=�	$aC�t��$�&�7 ��T�27b��8�k#�[�����<l��t��A6K�Q��(��@}d?1�2J��V��*M3ë��;p)b�W�"���5�#nw����uT�8B+^(q��S��Xʱjrۜ�������[��� y�����>�H+_%I<��0�^�Q���Ƹ"�|���-���GK7�����7�������f�*=�O!�v����#�@��DO�Ov�����Eg�q���nL5��� 2}	��W󾍂c�3�V!�� �4z��Y�����H���яH��f� ��,辦�jt���8jp:J�A/u�,ߒs��bz{��C��Tߴ9gd��� 36�gdH�%����M����sJ(>��9g1���)�RiF���RbO�Q�֛X�ؚ���}:8p&w���m���p�-����!l�0��Y���3�"�$ʱa��k�^ѷs��j��u���	�Q��l�&%�'�v+kf3��;����e�`,�ņ�}n��F�q�uh��Fxk_ ���<�$����p�0@�љd��*�E(��<殴ZCX���GCF9w5͸z��" ��}�����V`�b�0��y���|/���>1˦�Spr���w�0Ɂ�m��8{̔���>FT��L7q��WQB����
��,���˹�TRT��!q��
@_��W6.s'^�;݅0�_����̅A�,n��#���ѺV2h^Sw'	�,$u_���)��s���/�śg:���(�-��lg�o�eLp���j���Z�DG���˼p8�4��D|���`�-�>�|Ԥ�庙"�	�*0���]o5��,k7z2'�-#�����0��t̫�y0��x�7Jo��Q�:�AƷ~��$Q������	���,rÝc6r)���I�qw�������y�SyTN�_�G�8�|��b��uw;��G)Ȍ92E�6�3)����=/gfE�O�&�A���uD;�mat[���T�o���z��@#�V�'��PYِ��~4��g�[�����kFU�{P�J;�����Wa��^�����e"ǡ� @�M�b|W�+����dہ�RQ1(`�6�F�Lw���~�T���q��a�r���@�*o�0�'���LE�Q��n(:7*RE�;3'V�@��q��S@(aL"��q������ر���[qF�*�2�;W�l&C,VXj��2 ���7�O��G_	�gK$u�� �d��R�����x-ʿꦛZ޼���Q��#�o���s���3[V��\�;;&\Ln���Y�}}�X�D�.�ϺF��v�Z>'�1��M�\5���ER.wt�dֿ_�,z��=S�Y�h��;��z�М���AO	A5�z��Y�Ǥ� � ��ę�ZOv՜<��1W����#Y_�:��נ�O.dh�����+-Ēs�xZ%$*����s[l������;���)��n��
�If����{���6�Lt�z+�<)��u12!j�
��f(��*x3/�D6���Ir�L�<+.^	th�o`&�����Q�6` C&�A��:�z�g]���U !�D_D[B�6yЪ�g�#�g��\`�7f-q�ҳ���*:��H��Q[d1�g�*�yTֵ���V>\h4�h��-�sP��hd�kt���oI�>i��ȶ~�T	nZν3�O�2��K�&�_*��8`��W�� �Lj�h��
�Q�'�~(�;���K'J̡C��h;�,�=���.���슑�˨1�`J�Ĉv4F�7�	8{�-�ŋ��&J�(����N^I4����b�V�A�k�>�Fc��*�9�� r�A���1q�Q�i?��������2�">ѐXF�B�h�~0x�~���Vw)���9�2B]rv�=�T�˒�6A� "m��o��?���� ;ş1���g����Vj-�n
^JPE�i�$�o���jړ�Hr�Q��Z48�kb��K8�^��8.A��T!�h�|�T���ku}�..4�uK�#�j���~PIд\�+s��n�ֲRP����R�[�T�d�OJB���g�i	K\��l�i�I\�s�W�S~ʅ(��Hm?si�ȋ��dy����n�,��?�9W�K���o����ޔ����Q�($6i�w�������x���I,��<�>���c
lL���v��;ҫ��!/��X<=���#���0�Y�Oް>y��	oQ�a�Ӯ_%� �@�ؚΩ���בEXe\k�Me��w���v�i�3-;T�Q#�����]g͝�Xxh���k��O�!��")#Q;@ ��(�
D�x�	��,���s�j���i��U�V��"E�x�G�`��M]w-��K��`|�F�3{�>4������D�e�/�nү����}MC�gh�oM�E�E��*���U�(����4��,p��i��c��5�ɗ����bR��B�0��|��D�X�+������!|��:��`�M���0Y
�c<g&9��ύu-���p6V�Ѷ%sJW۷����}��+���n�bR�$�P�M��S���Vܠ��s�`��o{�¿�y��iu"[�ӻ��W�8B��+��h}b.,L�.m�W:p��xҊwn!�	Q?��6�q)\1��\!#ۅʐ�� ��n%���P���ک@�p g�%��I���%�����R�����/�um��s
%��e��o{��0�DݪCev�
)�����W)qݻ;���)�Y'l�0�ԇ�^Կ��=���5��:3�2Ҩ������3*�W</�8��j}"��@�A�
wi唚��t����q2}��AD�~�8ILc���Ȅ�ͣ��( ��)&����[/��ε�P���<W3��Y�Y�vm���b�afF���䋷wW�ui�
�'����L窋J7��'�z.zR!֋S�L�n�ȭ�ՌP�o)t�sgދ3}��u~�"�c	jʩ	��;�f�}�C�d�s���ϯI:�v�:���Hb5=3��t�K��Y1O_�tI�Ǻ�%��
o���u(~U��N�����qx��.�i��8�Lo�1P�n��	l�D��<\�<���ie�l���Q&Y�ξ��2�Q��X�|(1s���]\�bF͐&bjVbj(K	V�	�q�쳥ޡG�C8S�@F��(C�s�����K-����5��s��k
6P+�QK��/3Dd� [qoE�{��Sb��P	a�/a����*�M�$ �!j�[���{2��he��x�h�yw=DMtHë'��Y:7�$<��,��X����׋������ż��1���(��f|�ю��t^��_���&0 ��a����")S0�n�&-���Fز$@oE�]VAKߨ����(��pv_{�,���!�ݙD�Nh�������xH��3��Q�)�x�RW�V������1�#Y�29�,ee[Sr�1���,�{CƤ��ɾgF��J�Iɯ��@iF��M��dRu�{�m{XQw���&��S�#��3�&��3
�3����b�{��S�<��L_���4�+�wOL�����-C �b4/hJu#��S�{:��ac�J+i����/�3���T�8���:_U�3����o��CIJ*KHh�)�/fQ��O7vƂk��weЇ:�?�۰��Kn
u�%}��Y���ZxL_Y����Ǎ����S�Y|�6 m�é�vk���=���ۭ^.�C"S쭚��l�3�[	�@ھ�9�� �~�����F����Y��T%�$R-�2ʳ?�P�~���ǐ5C]�׀>�>/e�����q��ib����9��O�䐾c���͈�tm���UF��"��cQ��D3
�QB�=�g�_�~�ղf�9�)ׂ�.�?qln��YZ�ڙ��M��+���4Jh��!i���A{�=�������1e�
�%#,��%X~*�t���͐;a��?��t��û�_mxi<��4<����I`e��]AIB�1j�:wR'E;$�>tT>�΢>0�a�O�b�ݝ'�:d�Q�EQ��uݟ�RD)nxҠ�������ߞJN]{0��< ��E;B�]3!ܙ"��*���v��g����o4�����Pf�s3#�C�p�oa
}J�09�_�m՛Q��� ���)�Oc	�4��+��p���m5���
�6;���ldgoi���JgQ;���S 9��"�f�^T�yE�̿v�;����`��6�.��d�^ϼ���[�n=G#޵pa~��u�ކ���s������kI�9��g,
t,��Y^�Sۚ�ᤈ��E�c���=������E�P#��堪s��6�a��~ �'?�Ud�R��H��`eg4�[�S7B���D�Gg�(0@դ��mI�����YL��to$o��{������hKʻ?��Yg'ɤ��Avc��J2ia���=�m��CJ��MynT�hyI����䌙-����ǹ�����?Q����̨�+�?6�����s�P>���C��J;�'�ho��a4��T'�t>�[_V"nQ���mc���ab򭍺�Q�f�!���[���)}2��UM�ImS}��f�Fj��~Wj��'��J�v�9���:���TQk!��;5���P�C�i�1�ug忺�i�	��$��r�6��v3���l�zx�]���ڷ�� Z3�\�����r ��I���-�MA��%�݅�Zi�����暈P��SVk�%�y���0�F3���p�F�"��rnbP�9hWO�:c������C�vBK�n�0ΩzN�34�H�g�ͻK�-<��c�o������#<�CQ޽����n
7�H�^~�zWU�X�`ܨI:p�H�{��Dx����;
��Yf�y� 9���׷U�����c���B��M"td=�:Ҁr���ת��;H�K���dR,e1^懠WR���%|��	��be	P��#��p��{ln��7)��#"E�����jT�����Q�o�MQ
(���u�QO����u^T͡���j��v'� �i�}z�>��/f��"�[���Eo<rp:>��)x�g�8<�/�T��H���1�Pz����g���Gͦ�:�C�WZ:,�?�:�dx����t�`�4N�{��4Z��Z,�^����&�.��"�W��qY>��� ��|�>�ۙ�oG�p0D��u2�*��s��/k��9i��W=4�Wo�\�������!(D=VbȎ�
��]��g��(�f���f���*�jbB��ٹ#��oê�&*V�>�dt\��4�=�'eY׺����)ܭ衣�x9�=J jˆ��?V��[��=�[��^��J� 1ԃ��f;��I���`�%�8�@'a���T�U���77�`��'���%˲��K��Z�F�C��5��YG��RY�۴N��U��Ë?��K3�n�iؗ���� [
��H�K��Y��/ҤoM���"f�y�p���d,&h\?�G����2���aHuk�P;���L��b��+ۓ�3R6�S��)w��D Ð]��[f�Z�݉�ɳT��S��2���&nxad�{�HU.���畄"��b(a��¹�>�M���Ӏ���o'&I-�G)Uc0RWx�D�k�B
�7w��[�����]_w�$�=+(�8J�(�����v�p	u�i�*�~���np-�B���ޒ�#���\��+4Z���R�	��.�5��x�JoRkۜԽi�^zc��*#z��$Z6�������L�M�>�{Lt�J\��$Yټ��i�rn$*�c�b�M+�-Z"�*��ãz3���M�����A�+�$�+O`F�@ٌ�I�Q���ף:�a-a�����i����sm).k$��3Eڣt�P��G�=����n1M�~0�[.h��K�P�8w"@��(ܰ������g�L�~�O�bK
�z X����FV;� ��]K�wi/��c���n�ꈋF�$���Z �����1��-�.T��.������u�v�hJv�9����rGuvn�B�{���G��=AL���ãqd���Q�!P����̀&��uN+V"A�2��8`��
��.�I��{l1�����D�mK�`��LæS4@$4,����k�����?/q�U�H�wy(@)A鞗��	��@�i��q�y��$�;��pe��f��X��E"� ����k�vp� �F0�t�V�.���P��2*3�O�DqI����}�3n��g���A���i��}��+�N?@#� �x�]"0��V>瘺B���7D���g���lĈ��X��Jl�V*n�`$ۥ��@�u8�4�[����@��{�������}�L�V\�K�BE	 ����� ��$�[�1b�:̇�#���%�H�u*|���赵T���(G��|)/�m6���m�[�$��W�ⓠbe�E�P���x�WRMiD�5��wS�(�@K�h~by,B����Msm��C��5�>�+a��PܳJ<���n0�J Q˝)*��=�� �9���I�X�iO=Lgk�a�Jg���
�'�EI��r��.�#-�C����"�a_�||���$��Q�!��M��3�I��QaU=??�-8v��CU��A8\h��*-�����q���ӗ7�!�Һ��Ħ�\ϲB���
�$�b�񊽏Η��<�L'J[Ɉ���99�ODAԓϤӔJak9&�m�%6�P�o����tْ��qd B��P0���8l��p�=�=��@RN�(ְ���� 0/�0k�͡�0A��d��e�dv�M�8y������4��5���d<]4x���9��!���a�cZV�*��0�<m�W�zĩ��ȁuԭ�4��	\�c�S����J���]?WV�3�^/��z\�SH
�>�UVUvU`����\���n�0��@ђu��=g���*Z��ֹ�V;T53h�JH�wBI�zJV�p�"d�W���?�}�N�k�@�-�]�({� �_>pT� $�G�DF����Z���������MN�s�.�J�+&"9�m���*�B6�i�/Oͨ�F���-}����c%q���%�����L�q_�����[�*gFt�C���;�����>B�v��(�����_p�(ʁ�8�,\?0���y#��-(��[���	�Y]ؼJP�+yh,?$h�@�?\�n/�S�OV���e�u�S��*��M�X�uPe";o.�iTefsG��7?�;n�<Jr�n�-��R��Y�$}t��3TO����M�lY/�5]�����lVI���~l�(�5� z2�Lm��+Ss2$7���i�91D�(|��ݛ���s�80�[bam_�nlؿ8 ��-��5����~����Б����:/JE��v�q�8O-������[;��?t �w��!�
;�^�f{�p�F0]e���b�og։J[ _�ȼ>=�]�X������oMu��#�
���GL�I�L�����|Up2n���G	8Fp$
����E�[�;L�y�[ ��e��kcP���L=�^�e0�o9(}��FoQ#)s�h[�&#&�R	���W�#���h{%T|�h����(f�}�߯��
�$���oĄ��.��c�aL��K���B���E���Q��)$�i*���8'gW_KE����;
=DUңtAw��˰W�t��Z�i��l��.�_����KI��X�ѭo�o[:4%
�w���\ǩIc�<���Sc��y�w��>��Ҵ�j�N��w/w'?�m�d��$���\�qg�����u&Rv��p�-� uVp��d�u@^� �����+��-s@�R"5i���,"��p�P�X�&���uA��=	>�nRG`�&JK��_�gTS7�&�)/��["]����=��pn��^hUt�$$�TRb��A������������Y[M$��H!��QZ�L��gj�/��(بxAi!J�>vb�nn���k���,hS�������N�৒
,�s�dʠ����@W���V����k�
�<W"~4u��.�@st��� �xe� �R`'d��ÍN�g��<�h�dE)!�n�^(�a ���!�ۀ�~p�pyص2�'L��㙥���{�$'!"��L��f�U���RN���B��p6��b��"g��mge�{	���H�j�`!�\����6{��$T���sc�×��_�P2&j��)!���>K
�A�C �,�՚+�^U^�% ��o������K��Q�΅��"<2�$	�(,=��V2X���10���c�M�>9�S���"�<��b���n�a�;�ŷގ�X�ͧ�7��=�牳.i��5�~�rO٦��2G�_fY";��Rc�4��=CH����1|*):[��P�
��/�m��v���O77��'��bb���8��KӒ�B�t���3�%%���8���E��-{[m�;�i�BlkhҼ�6�i��"���B�Zs�&�C�9�8]��c��m���;���u����;h)8њe��'D���b��j��@K�ȃ"��n����yƲ��k�^�V�X�`.8��=��,��q�$�A�1�;7�dFwCe�|��{יYK�@q����)�写h�g}�PP���Ո���� �
`5|�t�@q;�WW�7�~L^�$ϔ.:$�X���|X�%���YT\,��`�Ys�f��I~������@��"/��A�����쩹�S*�(ۡ��'a��ۃ���y�;�8��;�C��<�
�A��E��θ�'�?�˾���S���Od�����w�ٟ��lA|�^� ��5��Ӟ|�%��Y����)�U��������H�~���/�gI�Y�0\'�%n����|o^��=qIK�##�d�D���C!�
i�;K��[O!�����۫�^�S͒0����H@m#k�?yo��0���2m�򓿣�����'[��iB"'6�$9p:e��@�#�݉��Ul���\�۾�h��k#E�VTj/K1�E���}��*���ǘ]�X��U��{ښ����Sףɨ��a.ߗP9t:�+f� J�6ܜ9]T�]�{�aA>�ڢ7e�/�F�'i6�y�/~���=��b(d�
��l8�6[q��Y6�^%����j{��	_��<2�h�7Cbb-���hM�lE���jy����6R��Yg���
qA���=�߼��;F��j�~�h:A�.â��sB+�pp�/�R0��V(�h7��N��N:�=Ļ��M�"�X�s��N�{R��BƳ��?A���f$}�u�1=� R!߀)���]��mB&9�����ՈڌK�C}������(Z3[��^�]��ԏu��~|���_�J����3���+�&�XO��W{W'��"�+�$�S"�s̤r
�A��~�@O�r� l��9�,.�'�G�V�ڦ��0"�e
�`z��z��ĺb�b��Ƃ+���vB4Ɛ����;�x� &ߏ��y�K�Y�ܟk������ĕ#��G�Kz�o�{r-s��($�3 Z5�ErKZ8��(������6�~�� �e���L�&�2ߘ=I_>-^Wd�"@q�*�4��������\6n.���S�Y�@��Dɩ%p��'��L�����bJ���af,�P�au�A�Ĭ%!���u���8��!Ыj�[E�QPqf�S�>�)��ީ\�����;-��
��|Oe8�=��Ҁ��^��Y�|m�h.���V��IkbA�����d�{�w��keQ�=����������fo���7�v!��ڟ^�(�޳Ĕ~�u��_ͮ4: C6n!2P1X;��g�Y$�����=0�T<7l�0��[#��$_X��	���C�����`��()8��2d&��iv^���!��=�9)n$�t7�/�:�ւ�-�\���l�Â���W�8[Z��g��Q���=Z�pU��Px���
'k)�5���C /H���V�DR�$�3������� Ddc��Bj�����W�}s`÷`W�g�ǧ*8)iJ�"a�^�ѵ:h��ڙ Yꉠ�n�_�5�n�G�A+�ը�?�e��bB�L$�k�������ޑ:���jE��~a��9'��p=���ۓJ��4�\����{`�i`)hG�mط	�%�Kf�� ĥJԬ+�}�P�f�[�0Y�Jp���,*���Y��/3�}x��8�������Jx��)�˒�{���QOƣР]�j����<J�A}��-�Va1E�3+s4͒_��?����=�֦� g����{���yyw�����92����m+��v8.�d�$Ł�6�?}���pfc27���h�sr���ޡA¤�3��A�]=J2�j�7�ه=I8;��I�ne�����#��ȹ�)QN�P�t?�跸~���-#���!?'_ŋ?l�%}py~��
����oH�h/���C��.
�y���/��j��	P�H��ٹh�BV���;qs�8v2�eAyrϣM���5��NA��B�Cܛ�?*���>�#�k2�R|������-a���Ѱ�ƈ��z֢1u�r�u�W��F]97�7wu���U���е��Za�u#<8S̅/D������l�������O���a����E�q�o�
������zN�^_�����Z��fa}�t�7�t�"O�}`�U����E�3|�Eם��$�˒ʌO�e��p1uW?9N��w�%%y�&|����E|�QTƚ��I̘�w�e��J��U�jv�oRV�B���Z���w�	k-��A.޼�Qb*ؙ�kJ2�3�t*�c�5�'/�'�̰'ջ���;��ª�$�����8�#G�W"����Hu����7��O��X��&]�Ի��)@�7 ���w�P^WM�)r%gT�*��'z���#.��I�N�?&�ڒ���t��UR�0g)T��(g�}���n�br�Hu����;٤�Tj�[���J� ��
�`��B�B��pI����n�u�|'RK��`23v�V�����	��<9�|�݄��u�K/䰚���n���v[:`�&*+��M��b�[��c��C
?�bGq��WD;I�:}��`8�7j�|�P���sk��8�q8��A6�ǀ�M����?z�"l��ޞ_+;�gk6֢�7���������-DM���Kő����It�H;���į
A���1����d�ՆǸŵq�ztG�v�Y%z����\e�Lhi{1>�98����ua򼢈����V�!�I|�hw�҃���H0F�L����HKs��EwJ!=�uk�E�>",����6���>�iq��Ѭ[jM�,{E`����!�)%עb9���r�UuX�>F�Rg�S&M��EK���6f�� �?� �5���!zX�`�:��_r�~�Y��j[|���Ab�گ���2Gi~A��`����I*�O��P�@��4y�Z�p�۵X*�|��D�ZZ��v�����zܿ뚱�c�e�l>��'���)�����C�?��g��-FE��t%���J �� l�J�U��P:e�tIA}�u�K��`<f�f�8ϖ@�^��
J�����+m�n����@�$/L%�c�������V�^Asם�A�<@ema�(�4���$��9s�2h�5��h��ʶ�ч��	{ٽ-f�'�u���]D�}.����i��tc�-\�ܥm�r�ƀN �#<.�NL��&�~d�+Z�5��c麨�� �r�4�Y&����*�6h(��WQ�#(���<A��O�Zơ*eB��Ts.�0j����D� VK�3���2��:�g�p��zx��i�Fr��==���|'A��"���n
d~s�K�	1r��ɓ
������_L���)�$�~�ufo\yv�}�Z=k�O��<�	>���M{��j1p���e�+��'-�N
=g��~�_ 	��������,bY���'G�\��2]�`d�p�	s� ����:��H"�J&�3w���γH�X%�/��Rߎ+Z�
IJ=��+���h�C�����'	v���)����<$|Vĕ�z�,��%e�
��������	��z���&mČ1ϭ�]�/+��ޚƶ�1/��_�^2�ʟ¬x/P�������Ƽc�xqyD��ɱ<��l_��M� F�ջޭg��M�9}�����N��dM�_nԢ�H0���=�uG(��m�"�W��;
}ȩ'�5$���@KF9(%��
I̊��x�޸���zl�O\J#]Ҹ�"j��J&����Q<��rW��ak��+49��t�?pސ6�|���0	˱�X��@)���#�6�R\�m��Q�%d�y�gC���
������v�w=�"����<����^�cy奈;��g�S���M %�N��b�ݍ�����U�5õ�n�s��?�&jY�����?sGq���=���Ol7w�(�s�� |b������l�9�*V�K�dSf��&��{џ���g�٤ky�՘Hߓ��[���؝��	Q��<n�\l�+B2��2�8(���3x����im���:�U}\�D��͝�zb*ss֖���9*���?5u٦�by�ZטA/���������;�Iifpj-DfM�[�U2*W+� ��1,:�k>~��?�ئ�PA�T�0� ��~����ux������8�W����b����A���K1�2?�������W��R�)�`����4�jҧ�4B�X�@�H�@��B2��,��}�G>��(�;�n9�H�Os�R�ѳ�{u;��U��!-7��H��i�so�6������ފ���Z?G��5�li��6/;��.m� 1e�z���T,}�n5k��)C2�?Ť/�p@�v�RghO0���uhF~f��N��mo���K�`g���߾���-\y����J�G������y-��钅3�L�_Fi�R0�q���r�!~�u(h�ys�Wq���}���3{����`\�d���I�͏��ʘ-��x�$l¨ܽ�|sz�:�)�K�W�B�����3�e�/�A<c⶙q�˃EX��W��'�9�0/2�RF�V����{��Lg�t�b��&f�æ�j�%�G4ΈE|n�9XcP:�`���!���.�ea�3v�x[KW����_�1@�	=3�l�IV��sd0�W�ѷת��	�c$5ށ]����F���$�h)c�-$�B)4
�L1=�߳��nƺ��D��H(-�zo���pt�	��{j�[��D��L�9�>Q�o+�*1���(�Ur�����^K�$�#���֪����=OK�gT��m#@ָ��B�|�����!��&u�ʆ_�Ȗ/�6������NN����Z�	{�³9@��<;�FWd�M�� �����9.u� �cs���g��{�}0H�+�u.����T{.d��	.�~,���Ǟ� a|8���>z7^��)+�~}�g~X��zKx��1A{�\�ك�<|J�9��(�����ˑi�8_�-�����z���������s�w���(��&a �K�h��l�	�H�`���d�
^p1(uz�XS�8%}V����0�h�*{�`'�|�i��Hq�S;O��cٱݝ���u��0�~lhs��&	�����\�l�]�f���ϔ>������7kr>�\��2B�s��4�2!EB�͞�9J���)� �}�:">�5� T��F,�@��D+��KN��d Lm�3��2Ը�ϖY�O��s�����z&�b`6Q)���A�������=��w��u��,��9��DNLz���L�<�'���Js]W��'Z�g�AS�"	a[:.�|�BvV�)�Yq��`_Z�W�
C?9��kv�=�3���a�&��2B.�,!���؀�+z�فI�(�a��gh��=W`��$k��*���ak��
(��c�&�qU�%���uwpp����Ϋ�SHG�hm������"tr.B�@�֒��(4U.h9S����$o~;�u�X�ai��:��E�	��\rd����P57KDs�ª���'h�����Ru�aj�w���A9L�ݮ�03�g��;1*6���ؔ��"�.��#��Q��=:��	���Ŝ�-5�������jgě��W3l3��~_�A���'�j�G���U�O�H.3§�
���m����i0�t��f�
���ݵ��U�QE��yT�| 
�
Z&��NTM*B�Y���

x?D�|�i!\H��E�;�Β#�0��X�"����s�"8\�~Wr�5�9W!�ш42���W!z��[٢���!�!���_�>H��'��x)���;��(baj����]���b�-p�}�<-Bj��3�6%�D@ڿ�q�\��w��E.���'0��ʥs'�NĹs�~�d[xr
U:��4?`�FM�ܩ�n�-�5�iG�s�5ɰ�6�W{U����S��}�P��F�<��C�e����dA��AT�ً�q��T|�lP�����a���x�p�޹��@<�z����8]SpP�B�P�;����k�!܍���E:�Y6^I�?�V��]��^�M�sN\�! *����^���0ō�׼V�b�Sh�J��'Js�7�?�Bw� �n�
�8jQ���,> d�J �L.�6��d�Q�H��&�������}�nLF����:��F+6��pD"�_�e	<�g�rjbk�v!����K��R�D&�����,*w��*�l6�H���Xri��[�O��Q��K��=�LV��<�=��m��CH�"�^c?v�/�=ˬ�|95IVԍ�����)��^�{�v]����$I6M����A��[j�41���y������)�Wsȧ���ݝ�{@̂�V7r�����M^ɹ#0VT�ɼ����������ay,��L��|d)�����?9�S���ߔ�nR[�Т�5^����p�N������Ү�8
T�5l��&����=Bk�y���N|��{�A(]���������J�Q��q���K��Ͷ2�/��@ŀ�T54����� �>��,��&v|@b�Su�Nk	���E�T������� �Rڮ��X�"����.������;T��V���^(�mb����9�i�>2�?L�F��C�DvS��;3kC��pY��>�֘������	9��44�X�_�w7�
2�M���5�)V	�7�S�e m(�ѳ��ɑ���9�������)r�Ae�swGZ�����Q&�A��9��u@Pp+�s�s��X"l�cS/hy�-�z��&�6wT�#�K�!i�o܀=�����h���&ơ_�PN������d�#�<s��b(n�~��	%%�!lU��`�ME�P�Yd���5L����vכ3P������S;玲�>b� ]|Me� ��X�ߌ�}bI����׶�>K��������>kf$��|`٧vJ��B�2��1 d
����U�70/�Q�⎚��2w!wI&�Ml���Z�$�t��͑,���EF�/�Y�3�����aJ���?�����-�`�xǧ,��"aY�$���N�b�(�!�d˩��_o!��D�aZ��@�K������K��w�2�׀����3�1���{Cg���k�/ ����xW�鄘��YՃ���c���V;�S^�fI͡�x�pW*pĵ������@H/<;��els<ҵ�M����8�
+b���\�n<,�]��$<e^Y��Ĉ��!���O|c�^�-��qk�Q*n���^1&C���§A��q�4>Bͦq���%VAx�Ӆ"���)��L���S�?�J���
O�Y��H�~���0���)ig���d�ǻ2Oc��te��\�����s���%G�g��.�l���u&��8Ѝ�Q֞(�[5��k[Bez�b]�^�!���}(\_��p��]�����⥢W���`���}���_{�e��z�Q�����v���޲��b)+��h1��*�8�R����Y�_?��.eH-Tt�4��)�%;�.tӓg)â��V.
:k��4��(3^�6�c���-~?j���k�� me�n�	c�ʬ���?�Ɂ�X+i���{;(;9�����I��7�����F��<H�D�������.��2+�%��>� Z1d=���A[�v$!Q�X��W�rJD��/�	<����?�^���M�����M�Z�r]��!R� ����)~K�ttGhy�󜋛�����������&�qG�u�}0�x��fՅd$��B3z���t-�I�s� T���cJ;pU���䊏yt9_J���Z�نHZ N ���l�?,�',�DuS Y��J7�p�[�3�N�a��F��FP�7l̙�U$r����Ł5�Y?B�8U���F�v��s���!�����_1W���ԣ�NЍ#����+T���8.ow���nK�4̺sӂ�8L�])um"<�G���ُC8��:�3����Z�m_��#f�0�~�Jh��<1<��!��9	[��N�֊�4���m��3�9VU����PK[��<��P9�L"<���:�k͸�}5�3k�(SrI�����r�r�漖�CP� �i�/C��rD�"O�b���0À�i3���T�8�OԹ�ꉮ�#s2���Q��yLX�9.��U�U���ubݻ�8������7j��i��t�~^8����7ۆ�Aii+�O�n�Ov4�AK�vY��T$ާ���X��k�Aٙư�g�h���o{��@(f�y������-��G��rH3{Fڤ#�?�V��=��i����6�C�y�E�!���_g|F�J�?�{�"�G3�T*����1@�a4:�7Ll���y��E���ɵ��~@:/�5�V1�$�q��;�0�r�&]���uʓ��d:N���h���1��|��0�'=:o]�)�r)i�8�4WC
4�-@��L6��V�LڮԐ0�VX�*a'�"��o�acj��DEʐ���\>{#����,	ao<���z��i����Cͼ`@�S���7={,yX�]<���S�^2�k;V��F]:�r1�ʬ�b/=y�JR��M;��Vۃ����?��0��vH�h΢�ڙn+%���U�sa7Zٚ�ҍ��~2n�p�Y�PA���dX������X�|����9�d�o(<W�67��s���5��%�����	.��	؃ì[��?�@�����1�D�1!m�5u�&�x���<G4�=i�ݍ�i~-w�P7Q2,l��Μ*ɓ����t��|��"d��F��J[��?��٢���8���_�)G���L��O�� ,Q��+n�$)l6�rd뽣�i���"�f�K��K�{�M�ݪ�q�R�A�}���ϫ�Ӡ��*�,���_`��(�j�3B�{���J��*B<=lr��ydȂ�p���[�Q�Z�͂'���6��~�×s�	���ݓ��l#���W����pNDϮ�g� uO���s��T�|�6�y:e!m����N�ϙ���8�ݰS}�7~U��QGֆW�LɃ�{t5�FNr<�����.N�X���6W��K��UL���5��nfvmgG�,;%quw̩���'�Ο_�)�IA� �+�2�W`�����T�hn��?��Y\�lX1V�W
'=�ܙ~�'��0#��=���ۢI��|�k��RQ�P� ��0�W|�
l~+>�u-��Y�>�&�p��B́90����\���q��j�+ �q�JY�� &�Դ�ulK����^�0Ӻ��o���G=U�CI��G�y�y�jS@�������#�B��U�y�Ѹ�{�ZlE]x4�	ԣp�B��FI��1��SU���l��Ơ�|,��Af��o�IX{84"�ݢz��� ����i2���[Z5-o�<ɥ�SF�Xn����@Ćr�?��D?��U�&�7k�o����q�%�[ �5K�[$�N�b����O�aE^�r�+Ah��MX���r��N���&l�"}�.��"���E��7����]�82�--�6{��UQC���Z� Hs�r� zXh��b����ĳV����<��#]���s��!�?�F[6ǯ����c鑒p�*���5����gP+�v�����9B|7�Ƶ��@��qۤ�7^8����������2�#RB���Z3��{�Ӭ~�vg��o�_����t!_�S���d�#�������>�),�ȶqy�:d^�9�rGGU�� �K�K����~F�}���Jʟ����<�im!�?6Z\�%1��foaKQ��֔'�'���}k#��z�O�Pn1��[|�1��=&;U��|�Xu)�>��j�
m�Mn8�*����m<w������&­r�ꢼ���J�V����0�2����IK��O�>(k=��Qy+$-��#I�q�g�a�ygD�t��Z��"��Y���>Y
��D`i� �v���DHц��@r�Qg$��J�Xm��&j��M������ΉW���Z��z0ͧ�Ԧgᐲ�������o�IS�s�_����#Vm/m�>�%`j#S�;�!���A��όe)p\3��rX���9��3'���IPx8�v��tWX���U��ו����&@ȗ�ŕ>���]YG��a1���N�.�����x	YW�-zM�t�v
Xh�d�5?��0���H���`�$`0 C�.�m��r�
�O<�ê����|�rHJ1!����O���Ķ�W�PT\����(�v5��������Nٿ�� RRB?������=��P16�}b �ԛ�U�1ð�k�!>��� 3�bD���S@�o�#$덏�&�?��A/��]�M���v���_c��ԅhH*���ˑ�}׉��?�q#(ܿ���N������Kund}9XgK��z���~�#�} � ��ϙH�I6T��A�UP?���I\ZD�ճ��S'�6f&]�y��a=Z!+�)��K�{�Y�\ol�tq4���!�:�db�;`�,N�*�I��cv�(q���aQ.@�݁���'+S�s�*T�����<�mR�5wX<ǳ�F{P(xn���"0�n��ϐ��!e\f�mV�h��,�e����m�n�	��w�UATųf�dtϾ���y��y���A#[�pα������_׬� �~��X�p�.�P��gTu`�'�\�]�viw�h#���7��-z���g�l�fD!�w�lr��!��n*<ۈߊ'3�J�
ǝ�t��Jk�$����pb)A�U��|�E���1P5@�(�+L+L�+-�S�&+
�\� C�����0�~xF�4��
�#@Y��������m8ĝ�Z��/��� �]M?{��/�!�VLʠa�
��NX�W�y@Z%E<^�<,�����mvZ����� mh�18j>���f]1C{���'�Gw�(`A�l�K��Q���`o�k�f��w�(���2
����A��U�/�wy�r7�[[!z��:���۠��)������yj�K���O����E�@"#E�j뵔��%��Q{��&-8{�f��F�~AGpa��&Sb<"��q��|Uu\�$��0�}aYm�+ P��2�0���y�[�h�@h��nk�I�}u7����@ Od�&��o���e4��vcٻ��-#g�:�~,���Lf�D������πr7���j �5-jx!QS0��#Hy�$���bM]�SQ#S���z���P�����&e���$y�O���RסDC\X��ʭ�2�r��=<�]D��ge�IN�f/�7tO�O�I�߂�щĥ:�������S�L���q���{i��:�vl�jk���wRS���s~o�S"윿nӽ[=��;9.��	��	k*�~є�a��*
��P7�Y4!���[�,ټ�3%�_�Q�f�ƞ��rC�s���M���nU�<5�P��S�L'(��b�J��/O!�_a����U�����>T���֟�Ճ�e=��CB	l��!��q��%��n����A+���sA/"��@��@���� ��R�s����K"غ��K�߅O���P�5?�,�U7ߚPy2�GR��>#%7�YHЮ���P�#�)HN�5�x�y~8��<��zo�öZ1muw�,e1xt����d8��$�ʻ;R^�V��i6l ?[O12<��?�n�h���n�s��U^ɡ�z}�<H���{^&t����7�KeN�gL	� �O֜$wU������pBrp����3 ���,7M@��ܼ�࿔cE�2���e-�P��'ݾ� �?Eҭ�`�c��}|=�b������B@=j����<�-OxfDOI4�Hc>G!�	��8.j� 'T�@�C�:���(�N�I1�C;  C�^k�%<Z���^��[\�/Q���B 5Փ�Q�W{Lwb^�/�9b������<��i�}2��2-�+�=2%�@F���Sb3�
���' �&��1\F�q�l��C���NS�6�G��D�m�W����9�l9e9��kA��T�p����u�;Q��~����>F�vi�r�.�vϣ��<��#��x�l���)�F'�e�~�[bl��(��2w�/ސ堋������θ��^5��h�k�������ȳ���������kx�w��WЎl�T�:���pe������g�i��K̏��[]#.�x˺K����(f�}0�G���Ud�5.e0e��z�G�������-�~��]}ł�e��F���/>۳�u�س����v�쵑�����[�:��js�`�\�S{!�'���#ψ�}���w��~�/�?����VlQ���?������lXzZʡ]~zڴm4P�J����1˳���.����U(�*��L�z�/V�3=�D�Z0ߤ/�K���!(�k��)t5�wȌ,���.��
&i&����?{w;���ࠅ��_?غ1y�
�s���X�.G��1��C�����YSc��/!.l�6��f��X�׮{۷< a���@-�u{uJN�iq��u��CP�	n(��cƢ�xkѫ q �N�^J��[� �\�\�X�������;���4�QA�0�����j����cBe�����G&����G���D�w��$�|i�Z��c����V"~!\��g;�Wol�I���X͠i�aa�*�Ĺ��+�Z( �����du91��A{�$�����N�˷�w����.#U�{�+?��y��Qa˥������"Kv7Wa������V���y��ש��+.��5�{�ζw�v6�Hh�-���%�CW#H�"%W��НIS+��j���ѥry��Y����hźZ���q��	p�L���s����2��J=Fn�����^�z0C�FH��CK��rȱ��S�t&)�aoE����ʂ?7V�#�TT<���v�}S<^I��zx�M"�%�R@����w� )���Ƽ�oދ٪S;;��@�n���BJbk> �4H��I��k�fa�H�m���Y2��YcD��!o*;h��\_���>_������9��nu��x�H��]H8៲�D���6w�����P�;����/r���ff�'����
�4�M�q���gf������7ј��Y~�U�x�4�1���c�*�/s�w�S]��gii�4ˎ�Lٺ��{�����I^�����<b�̓��{ti�*7�F;���F�OA�i�#<.�������;�L�ʜ��OR����i�e�w�����J��o���9�=���74gNE!Sb��p�
Ч��DG�"��w*
�����Ę���8r��\���I�7&���������_�,�G�K�3`��$��6�`�<�*u��$5�O�!1�kSv�]�DVF$�:��\�֏�%d��W�M����j(cS����M����Y/xBx�Ij��T��,D�"�^��R�=h&n�c�]��KB0H�EZ�0k�`�)D_&��6`�t���O9O�%�+�n���tR�S�q7_5�8�\�'�h��>έ
� ={Ѫ���"��Js��Y�%����`-�i��(:�w���V����B��N�ugc� G��FeJ
���qN�U�܊��	�c5W���[>��`���O�w'/S�a�B"�s9����$�H�f�`|�eR��Q?8򙓢d�S��_��Y�z�>f��~����)���p��^?��.n��@��Yn��Ո6-�����!:�H���=�Y������k���?���A��Ū$���� gA�"�$���{�5�2����s-�mq�u�B#a�('R�9���@����[��w��*c�q���;��z~�Er�T�[}���6g�Q:|T7�h��� 4���ecy1���h�^��jⷾN��+�_H���0km8��k`?%i���4kC���T�t�>b�����~3��/�Y�"�����	�ht�X���j
T���2�7�XKh��2`�����N�d����Xz��M|��Ĩh�Ԫ��e�Kԧ����8�k�bא�����1h����k4ӹ��@�N1L=g��L#7����/)�� b�O��[�{b@�\�SΠ6�p�%&��k�[z?���1�a�Х��&#����O��WJ�ڋ��P�Mw�-�sS�5���/�$x���F���{�'s<��H8|���w%�D��e�
�#�+�}a��2ɽ:5�K.g��5��g�J��������B���4��,���drN�H��<<
F�y'�I��n 0�	��(�4�{��(.v�0�3�$�->-�߰[^�cS7��F?�F��5wH��^@�ϙ�n߀yB��}�ӱ~�pV��2�%��y�6<����Qg`���C�F3���
���J��������/Wh��{S0S��e��lOh�BH��.W�̡P؟q�tjx{�T�L�Z���~��;	1���>B��T�;�2�v�T��7�s�˧�{�̀��Q�&*�r�dA{g:�֛t��}Dl��ո.�Mտ%y�s%�0���Ծ����M�
�(��pz�lnQ�_k%�ꥮ��R�KW�+0���׮\ROx(D"����x
ۮ�&%����C2���A<п��}���c']�~�.��?�G��D S�K�;%�Z��-7�.8���<�^��
B̩2��^��/�!���y��A����&wB�]�w�ye5�񅯓,���5��})��L���L�?��<���0iMt��S����F�p\S��p��Q�r���Ԏ�&"���
��so�T���_t�K�� �\6�䃣i�ه�T;�j3�@�%��6y8�bi��;P�V!�TOX��l-�A�v�
�GVФġ��vo�c*L��͓ܼ��9�2��CQ��weGU�<��9T;�5S$[�fMp8o�ebx�����*A�If�ā�	��4S��:�� TK)3| �~�[↎=g���*���5P�9��؞�z��/��N����3j�v�34/�oF�l�#�����������s�P����cpصno�k�Z|��^v˵
vh"�<]q�h>�����`��i��b��S�D U�����޼�|���r�>Є; H��;�JiL���������k0�h*���u&f�����G )��(`�9�C��v���΁� ����ŀ��@��l>=H���[8��A���9Q���"�y��8�|54��E�<�H% ^�鸣ɥ)7�Fܔ2T�9��8�~���/2��7O��-�`�z��S��]�@2񦿏Jڳ����$d!G����l����|V@���*#�n��A��#�`����mn�}Ÿ�Ҽ�Zp�'Bv��|P7lx��ۭ]Zf$ �s/(�i4b�T�.>�,�<�ys��ׅQ� �Zx��?��]��۟��E�z��F����*]��B�L-I��K��Z�f9�a�����5��Q���Otؙ�u�;׬/���ʒ=�=	1�w�us��C`V�	�?p�Y��k��!�6�b����~��٢�N�l6aN�
-�+` ��t��-:S͞��L9���WDa�B9s$[s0�Y#�iU�5�[�z�?6��8a�uM�<�_��j2p�
�h`��rdn�#��-��V�lnR�O�=��	����!�%^�(��)8��*�#Sn�v���g�-������=̗�\W�¨���$���>fW��L-_��g�6>)�3H�_�X��X�WU!��Z�U���(�M�Z��\�rvG��n8���>'fe��R���KB�Ӗ�	���a�L�͠�Q��=���b���8�q�Cp�_���I��Į�J���2��)�fC^F�d!����@�t'J\oŧ��V���W2>g�dd�z�򘬡A�} ۺ��n�V<�k���V�}��V|�<���Y"d���d��H	�9@B����ʥ~�D�Z��m1V)}R��m�(!s�7��j���U0�-c,�8�U���]��R�*p���.�m�ڀ!�~�M�Մzq|����D��/���s��0��FD���~K,�˯|����-h*:���)v��sS@�_�G� ���i�U�껵C��x���@��^c"�K���Ǳi��8�`��.��9�̕Pr�'����)T�Ҩ%���������~��V�JJ��wCB�ǶHٜRS���!��C3R<q�u�P����+f����\�s�t_3���F�pκX<�Ʀ�sՇ��5��v�d��Vh����D������a@|<��o���b���*`��T!�&T���&���ҏ�/���3���J2�(���{J�ʾr~ϗR8D�ʄ�5T痢�~J
�޸���h ���5���S�F�6�*3�������C��g}�t7M&�f0�&Ү�0�H�b������Z�]�t�Ek�yˍ�T"��(R0��@�z,����l��&R ��M� �0J�ފ �8;�0��-4CZq=�'=Ö��dښ���f����\�%D���<�U�4SzZB�O�W1��_�"���c'�v�/���OAgxe��!�B[�`��`Rc���ȳe�!W@t����ƺHM\������~1Y�|���ELԾABt����9�7I%^�OV���Z����"V ���vs�>Q�:R����"Q����Ӣ�m�� �m%*��싧�Q���@'�{j�h��U�&� ��e�9'�dTĮ���]��E7�YzZ�4	�t�Ym�iK��9�J���#ȋ��(ĮR��Jp�?�[G���ED����5��`�_��cW�����>��E�,B�O��MU��xTG0B�ucv,ߛ��莟Xw\�t���n:,k�t�5���2��KF����ПCR��.�����F�)�
����&5ί(Gg�-��ə�'f��f?Ud	6�c!���"M�I�5AY�:�����2L��TGa���2Z�?U	����PM�nػ=�5鱨A���x�5��!ecqV���T,9��6�6��m�ԯ�ZW*�������Ǯ�ށ�W�ah�YB�W[3�͢?¯�� P��*\�*�hA����q��S梊Z|&Z'HP�涖V�s�֑BٷɌ�`��v�	Hʛ,�2��9p �]�UF(�ރ����3_q9yb� �w`�t�	�������8N�D&�,�t�e�T�eQ��7���I؊��9�`D�L���qs�|"�ԤU�Ưg�R �Y����erc����F2��v��:�	%��)Z%������1�8v�b�z�v�s�#)/����BP�ǵ�Y��= buF�߆Ǒc,��(�/���g�'����#�Xg�^�|��/��O�A����F��D8N��Eoj]���Ћ�Ơ����f^z��x5��g"�9���	����B�ŬX�$;-=��-,~��L��f�|{�w��B��mh���@���J,	3 I��O4Ik�>��6a����0��;-�tMd��~*�z(�hU�Y�	�s_���c�c�����cv �7c�Me��sT���(R60_�\uNl���(������_)�9�pR��{� ~bV;(Q�ؤ����Y�b�u��v��;i�Y�.�:��P)����E�֠��#�r�He	�O%˪6?eV��'�8?v����_�O`�_FBk>��h��W-��B"�Z�֟۷�c\����� �2uw�>><�k`���Ϳ�YU_���N{��P�BJ����q�N!�qCHyB D(c�����#��O�d���-�
}�_l(�L�U�J�`�6BO)}
wiЦH�нF��T�U=��S�>����ێb��댡�^��8�ñ8bW�~x.��0e���D�)(���6E�'�����θP��b�
��iҌ��G���/4�xK��c��R�k]�����;��q�oa�T��B?4����l�ă�_�Iaː�H�������3�ne�JE�IIg�����S��1�~ 7Y�Y���ī�尣�18���λ�Oěw��٧Q^A~�l��r4ᜲ���
��AOch����˹Ο$��NIvO��� !����'[�+�86��F%���nq��4~�P���{�s�ص�3搒\]%���� �8�s�������l�hd5��l�����3��J�:��i���r5Uqx�!�����T��m��-����l� �F-\4H�NCB��H�:y��>��8�>�s�{Cݷ��G���S�����@q� A�1��O��(�c`��.�:��Ȣ��R8%�p��w���A���:i��[{�[/���iD�*�I�R���QY	Tܣc�j?�q��9�^�(�w:lɛ	qU�ݏ��B4��{65UOԾ�6oV�T����f����,â:��g���6�xZl0
/�V8ra����T2�b.jW5ɮu��t,
�	�m��%��5-S�/p�O�A8���m���g���� +�-}�?bޭN��g��1�o9�LYk��Q�̀W�hݖ�CtN� ��.�fu+;�������.�;N�L+���~w�����8V�|�l���:�@���j�\Q2Iith�'���tѲi����eS�)(��0#�-]��I)����^�T���:*���Ɨ�7׳l�0<�u\�D��r�Ŧ �]nv�&j"���}�� �+�,i����1T����2?q+f�(��\ԗ��<~��BnG)�
�����!�L��FD֔��\y�'�}0����Eq����L\h]|�B�J�^�<�ch^�ӓ�/��H��!	�CS>r�x�5<�N�O��p�vwو��L�x@��I��,��|�J_�:���A������3U&�A!��xF(���]�ȡ��CU�������:	�b:��\�g,Z��y�Z�%�~+4O�X�w7�N������D�%ZȽʡ����6��=VF7�*�[��ǁX�{�\t�@b��p����~^������o��w{�StUu.���h"���ݲ����$�tO�BPp�\!�ϖ�/��*#R4'?&�:�Vh��Ȥn�%Q��$!֦���[��(�l������C�o��������ց�'H��q�!���S���.e���VIa�	?�1��IskGJ�յo%]�x�a��R��(�de��/`�B��6�]�I��BH�U�Ų9)6�6S�[u*:�Ry�Uuqz�޿���=I�G�z�L`� (�$	�H�(m'퀗��W����q �t��I`�8�pG��A�x!��ϫ�@<߂�&}j��Q�GD<�����I���밵��/.���o��=�N���6�W\b'�=O�aj�:"�����@dy@�>xDx��q@e�y~ �:HKF�r���-L|I��lIy=c��i���3<�$f���T�2/�ej4�臚Հ�]��$��D��ՙ}�`@��!�(�0�wUm�����ra��.x��J�<�-+���ǽy��_I�|�0�jff��
�J�4���h�O�6	x���(k�� �4���چD߫�<fJ鑻zd��������Ir�j3���-47��oT�¼���;�ֽ;���Hƴ�8�vD�	5�8�E�����TMp�;���ǃ1��V(���� z5�p��ˤ�:�$1����~������=�SX9qt��r2 -2D��: �@��o䢋�f�0FT+�9����MF&U;���I������G��2��)��O��Z;�ļ�!��t{Z��F�ޗi�T}���Y��z9nA��y��)Ѥ��΂X8�>��T_k�D�_�k<�Q	~E��)��va��F $��,,���,�M��H��]�;�1} a����Y�p���"k �z�$h�Ԃ��
�4w��7�sw��w�a�Ҕd��D&A��K��A�/XE���m���m4J�Z��MJ=.�*�6�q~�����#��#��ڠL]S���k����;�+s4Z]��%����SL�\U)��/�【��=��^-��@�n�&B�K�>��8"�sܥ,�0��g���C���cn1]Ɗ����!�f�Y���6���������-Nh�
��bE���=�P����*�=;�Fx�ؾ�I�HW��H{O�	P���1�f�'Y"qן;�F���ř���8;D]�,O:PX��I=�C�0�t����dJ恿 �7���+���jޜ��B	��ak}�oۉ�Q�T��Z �o���Tk���=��1�8-����K�!bd*?+׭%%��4�4�	*�{�Av�gbƒə`���,���_=R��+��r Aw5]�7����[rz;
����ü �g���������nk���Y?l�Am>�ΦZ�?�>�?#��T9,JM-v�h��X�3��bKQ�>L��
�8�/�����z�{e����;�_Ă��&6S��M3�j$���Q�֩Y�k����Ć[hk
yI�#�QUB�t6~W�p{�je�M�S���ȭ����<����{H��"���{��j�8�s�MRR��7�.�g�Z.��;�������&ɠ7�r������s b�q_y�^�j���+�?��mnH��^�LA�C��f���H
��4o>U���c�6��ꡲky�0M$��ƵVC�r�r'����#�P���5�>%���Ly��9q�go�j|0��L�%z1��3��~�a��|��&�j�v������ )��+���><rqb�f+,�T�$o����:�ΐ�/���=ܦ�T=\I�|�ӱ��L���˻�^��t� i�x�=y��ur�;a�X�[\?�:u�bgt،F�'�rl_�ȹ|���%��,��1W���K畟��\�
���u3�ދ+��P�~�@�P|�ׂU�`Ƞ��	h¨��r{��{oc���|���[�A�ׄ0���+�`Ѭ\sOY��D������Ȏ�z�>��<��P��JϺ��(fTD'?u#���R
QO�xR��$���^��V>r�cB(��N!�<��A5�.����\΍4~�1Ϣ�X��w��k���k��I3��@��`�)V^*Z��S�o%%!�����P����e�;_�J@.;�7��]N4�b�YS�-�%��bԔs��t���T�I�<�).��Ѓ>�h�����ͨH�ۉI%��OL�Qo�� ���k&8_�1ڊ�e�v 4����[s�qU��|���6�m��>3Qe*i���h��o���J�:kr��R�k9���F�,渽��y9�?wa�do?���Lbp�~oIf:��]��ox��8��F,�4��~���Vn"KKY^|�.lU�|���c�9�²AF�+8����
��m�bR�V&Ls͐\j�/啌��V�:S����_��@��O(���3�,��\��DH�6)�F Ν���7���?Nԟ*8���`(���>����B{�#��C ��������|�-[
�cVx�$V��
����J�@K8�<��M�Y��+���ձ�4O�rCK��%d	wDD�pi��Tޞ�0o���30y�@#D�W �������|�͕(*0�(���A�cR�WP�NdBf��Aך��-�|#��~�tc��a��������������~1������]R�(Ƅ�/�M`2���5V�5�}s�������SN�cT	���ˮ�=Q����������j�\jO���~��(���ҩ��u0�4k�J��p�I����۸����Aߩ�EGHRѶ���C�C?�0F��H^������a`K��Lȋ��`> q��t(�Q�-��ϥ"t�>���1hS�hY���kL�X~�DK�Ϧ��ּ=��x��Ax� k(��9p���*Wr�y�}f�������Q�
�4ei%9m1?��?�{�&�9p�m�r��oa"͖en/�9�׷Ϩp��:�tM�lˉ��-��+�A[��F�3��q<��?a��@?�x�x#��oY*`�!s�p��wW���9�n���'I9fĄ��}^��AY�T�c8uu��Le��U��g��S%�1�zB���[RAF���\D/����^0���V+�X+X��&|��
���x�=�����|���|��Z.kj�n�Tܘ��X�nj�j5(��ҬΡ�3�w"td3���i�Ѭ
" 0�$҃�12����J^n/K#�F}��C{g���'�,�C5b�Wf<��1`��e2��[V��T�x�;�Dȗ�ҕ����^ߞ���P�%}��g={Xz���B]}ϊ�13
�r�Xf䛽]�p����~���6�Z�F_S�t�.'k_��5�ʿS��/%@2��~Y_8����Ȧ g�B�p���y]:�o�AQw��Ҏ]���1Q�}8@}���l��U.\-��6[�=~�}����w� Y��;ѣ���9�嗔%����	u��;� C���\�Դ�M<��2q����m|��UM��'O\+����'p�����%z���M�A�*gڦ��z�X��t�G)�Q��Ϧ�<�������3�F����vL<7g�����88���uW��my�QE�Ohʋ'��I��^�����1���}�x�t��1��v� p����c��*zܶ�Wұ5��3���2���Nq�'ߠNW|<�OKn����$޷I�he�|,��s����I	[���LѼ�S�'h��AЬ����+�]n�4;$�Pw��/���N�<�U��`(c�a�밬��['c���_��?�7#�,�)��,}/�r�
��۶'Z��0/�+��/�\M[h�H�&`�msf�`W���8�K*-H�;�!�C(�Y�̈��E?�������:�(����j���_�M$��a	De���~
��A��UB�r&�Q���|]�UxR�?��:�3���#)��M�D�5	a�7pM����#�G1��6�
i��!�V�OXS�k��{S0���ho,~ ���TM,��:�o�����څCxw:�z���Aѻ���"��MM!���̹�k𫀀�C��+Q���%�^9<�^r�7�����I��݃y�R��pI�����3	`�8i�D%n���m��Ɣ�CI���a���y3#��"I�M�v�����,��?u�hޚ7y}y�(?7F�/p�vmvLٔ���&�̠���m��b���!����h�k�T�%�VL����_�G�eK	��ǿJ3l��(��:N�X�k1�Z`!_� ~,�ԩ [�,�W�1�t�����Y\hA�#�A�H�����5�ͅ��U{{���Bl�Gt�T�6�*�	x��s nũA�������u}����x�dT[i �7��\;tP�1:��V+P�[�(�㧮mP���I�0��Uy�;��a:㿀��9`f�*O74WۙD뎋G}��Vu�y�d�ם����K���&��B[GY4P^H��[��ǫ<�Hó����K��if����80����Q�$���J�K;���/y��	��,X\^A��$�D�i{���K��
F�9���OHyA��ZZ֔M=��(`1Y4[>�V�F0�&4r/ˈ�� .C�����>=���3]�kEA�[rSOZT����[����|Y`���vP��� G�.`#o_�MS���Yw}�.+�ޠ�ALήL�����O��(�m��0�T��2�|����.�R�܍0���N�f�83c����h����F�R�WKuG�*��]%�rB���'MqЂ\[^g(X3%�"_�'sq]cyB�A��M�־>��_cc]M��G;O�!����q`�1J�"��z���\D�(��A໲�3��[�X'�0T@L���ïg��g�ϲR4Z��<�X)�9ƙ89<
S��Oo�z�Y۞�ݗ����C�W' ��:���-�Kxr��o�)/���&o���-�A�Nw�3�N`��&�i �,�ǘ>�}uӉ�+|
4��2������9�lɆz�a�C�ݻD��@�Ŝ�_������NK�@-	�xc{�$j������)e�f|*'��
n�qz����J�����|������ڈ>��')���;���l8���݉Ǜޑr�j&�<�g�~L�ځ�E� -�~�?gW���Fت��#��q�]�%#30Ft�=�U��;�/ą���k�y ���wf=��^f��Tk=G�ax)���FE<������~�꽝
E�̛G�c����:��� <��=�>��x5]�To�J����������+��A�����ih��*�����Uƒu�
#��q	5���W����\� Ia�Wo���`c���*�)��Ϯ.���:��r�>����G~�f@�!���^����N[_���M�=�X��#xB�)�����&ۖآz�4�/��{�io �#�aw<m�IP
�+w�a����m�^�ܭ���d����H���7)3� 0����,��ذ��W��l`��9k�EIv#����Ʊ\��o9��s2T�� k�IjwJ��� x;a/ r���[v]�x�T���x��EW�2����6?TH:���7:�c9�5�Ht;�o;�פ$�m	�j/��`5V���#�=Z��X[1bgsD��v��!��x %�Qԁ��{r%i��C�rи* .6D�Z���|R��qd*����eޮ�̱�@sw�I���_���z���D����y���x�+��0*��G�4L������w�֣��Uvfv���+2���|G��*�'2xxx����J<5(���p����÷5N.���蔅͊zgq��79)��d%kTn��Z��D�:��%"�A*��W�A��u�pX�M3K�t���;f��=.=�Ԡ��X����({�J�U� ��\�<7XT�pg<)��bs�T�z��?�
P�@�/����Z?�<	<�����?����N�iІ���4��D��%�!ɠ��������ZqGz���I(��p��[��`6T�)����(�����v]��E��� <3�)!:������Q��QUq�<Z%����3��� v�ɴ\UV��x�t[#�mߞ�� ��;�&��{���u����Ʃ���I�Q�d�w���m=G�Ҷ'�o�*���s��SC��_�����h�μ7k2�TN}X�N����g��@��d�3�K��
��\O��b��m��m�N�>��Ni���
��zjswjl:$����$AUL�[�3i��ج&��;o�d��x��/�g
?�#�;����K��_��҂�L{}~Wܦ3�Jٚ�5�X$7��#lk�kctT�>l�ߙ���(�ia�j ^P�+{�������$ ~_��,�Sb[p���p�&
��9��d�C�����E�<��a-�F����v�S���%�oI�Rg:�������k�L���{ ')�oq�~p�j.::{
��i���(��p�9g3����
�Z0���#9����<�0��-�ic�����S��� ��ޫ�(�]���|�֒�yĬOn�4T�-��o�Y�����^P9�I�@�����0<7c&��ɉe�}�U��$�$e�sF��?RߎV1s�#����{'�����R�����` o��8���G:�x 7H�(Y��(��.f�����v����v�͜��)�}C��N�zIX�<�8����;���t��/�o���|����N@�L�#��ќ-����nH]�
�=w���*��R/f�ܤ�o.��IĲNx�#mBa~�����q$:)�T�Yx�k~#"��H�	�V1��nu�Әo�$��eM�-waM��w~ ��`p��F�h���(JS�)
��z�£.�9a��f~t��W.�Le���@� k�����Tx5�)\��$��x8���@�YR#�����,���
�5q�X〰���Jgv6���'��������Itw�զk��f(��ZM��:�����.	�dr$�ox(����y��B�^�uT:��m�A� �N˹��8��Rgqͽn8W�P�ܽ��CC�����K���G@�p0�$nH[q9�q|�`p9(�!�=B��l�w���K���I7�]h���v���#�`�NgS���{���@ۢ�i��_���8�����ΦA�<��}v�<��$���s��e��qW�O�I��K�o�j��k�<EJ��`��!�@y��#� ��H/L]�{�{��f�����wK�=l�
#q��/ΐ�D��&�Z�:Y[e�I���/��}�+a�.�o �6� e��QV���Ҕ������w>z
] �Åj�b,���{h�^M�Y�����]#e��v_Fd�m�je�������a�c���݊��n���M	p�DY�C�`t�!�z��HBx�V�wG���t��%�W�S�ϻ]OB���6E�`��	��,�[w��L�,R����?�ۧ�d{�����z�����0j��ގ�Qz>�N����Yrbx�۪,�S�f��eS���C&9h72s���(�*
*�=@$���=~�k�<'�=3�+��C�&w���̓��1��#��͉���6B5�������%����Е3~>m�H�x c�3�|LP��1n�@�_��I�'�K;��I9�y�zlp=lY����+��uR�����?�ܟ�M�ߧ~9�+�1T�����T��ըߐ���yͯ�y�F5��$ �k܋1j��+�I�R�$B�A��s��I��!'����`���]�	�qlW�������u>O+I������f �u�"��Q���O�&��tjE"b�#�@��c��T([����l�Q̓hH@�;);~`��q$�M�-lf-f�B��W�����"f�����mO�;����
�H��/��W�����X��uO�wv����N�D�"ة�֩~*��ʡ���;=:�!����g��"���e5(�xU����tr\q�`��B��/C���6}�&$��䜅����'p�ޔE��!�r1C�
��w���N;���P%Q�i�r^�)Lj���|�,4�� ���z���([�l��F=r}���r�ǽ�"K�#��$�����P�5�Y� b ����c�s���ȥ�r�ʸ�/�L�	[7�.�,��t�	7�Ϫ�qu�<ӯ�+�D����:��,̬1cgA�ri
�~��XKB�Z�E�0�s�)?ǹD>ȭ{�?\����=NOђm܉�]K�7�b�|����� [b4�����w�ߓ���2���se���i�V��Mob55����GJw��Q��q%ą����YDi(5��˷�H*�>�w�Jd���a.t+��ۆq�u��D�ܸ9��m<�h��4�c4��j�*�=���H��QxYAL�O���?�.���A�	��"�WI� VVQ�&I�vm�Q^0(�0�$�������B���#�To�/*펎��W��0���<)���x��|�}�B�{Mǰ�j&: 
�~
pp��K��.����~��1rH��Lq
��H��@�++XO�:P��El͏Zˆ�3 -���b)/��k� 1��4�S�V�S�fO2z�X�
P�E��w���o�_[�_��Sݜ3�V��-"�Xѕ�~�(��0âJ~v�����>^�4���l��&������S���܌d-TI����B*tk̋�w 3"�����.	\S���P	���/�R�\��f�'���E��.FXA���F��bd��o�Q$+�ײ� �F��$ ����1�����C��,{�"�sۏP�Hh�>V��r��J��hް���k*	Q�1�H�/�i�#��+GU�O��~��WB�-�������S˝x�5?Zl�1�ʄ�d	�at�����9��e3ܥ�U���,��,r*�2�['�'Cm�oU�?߫۰�u�1y�n'Sk��*��A��9F������Qb�g�z֚�HR֐ө�&�����.T�?��F:7�S-s�j);h�X�X��&�"~���R�8���=�P%�h�3��t�K7������Ă�b�~��m3�IW���W�h���܄���#�lÖ\Zp�	�Æ��� 
�7�H}0�T�N�*_��Ehx�V�9��Ri���/������}гv�p��:?r���QI��
�
�u;Xd�K�Kξ�BAY|?���Ewy.Q��l��e��O�vrh�U��fQX#��E���u>��yv]A�Z`.�� /ჇB�\/�yZz�+����%�lL�^3��)�<9fɤS�X��9#F����X��>�W�%� �w���~�OmLw���C��
͎P@|.ʂTY�! �O��ǮnW��X>���%Y����Z�|O#�����L��_����镇��BO�V�V��!�+�"�e	�i:�����ta�V��3��AIY!�"�9��zY�F�r�E���`��@�P.���*�}t.>%0��qb�A�,�X��)��������t����`K�ޫ�3��(�8+��������<YpaճF�#�im�3��ܹ�5�|�-q�~�JO���}&��2��V�y8�_G���z���� ��X�^� 2�#�Q��Ks�hP��e�xm�K铒:~���M[�ᑤM�օ������ř�ձ��a�0G���`J��?ؠEt�l�~�
-Xۜ�j�<��ރ0�?�fuw+���dx�2Yn9�{0O��o�����-�Qw�]Y�P'�"����iBR\�-.{$G��6x��( ���շ�k-W����f�	�ɟ�6�HHm��-���!�����D�r����KNg��H�1φ�\�@I�C��G:XAew\R���=��[�c����j�ݸE�q���"�4�^�:]��!�'My�1mԮ���3b�����&��`�JU�-�$�
hI?��z�#��E�(��!'C�1%ڒ=��d�-��)�)1%��"ΆT��q.:[�S_����kĺ*	_������#*���x纍��K8ʈb�S���)�}T���h]h�z��pN�$$��W�U���)ު�p;�Gf��ˠH�o������V�&����Z�s�q+:��xE��d��-� .�I�� �̱0���w�[����* �F�
z��%2�T�M/q���W����:Ӡt?�����Ĵ���v\}��^g�j=ր���Q~��B?��d2-�ܖ��׊�H��篋tҠ��Gy�����c m2��Wo>��`E{3�hJ����e�~�h2�s$}�������?�	-�ɳL<�k����%4O�9��`
�Z�C!t~?�F������Ï�`��O��h�?*]�1�Wf��q� ���y/DI�a	u�ER�f�,^6�oiK:�UG�4n���ul;��9�Ί�=�D>��bP�i�p�u�{Bc�'��u�6H;��=�6�:�'�%�5.:{i�V9���H�m���^�����<�)9/_����g�#�CF|��;�eAy-q�k�/�vN�����C[�K%�Rk! V5`���k��Jo����>����/. �X
���<o�'�$U���������j�N{%���H�
g+D��+�n��}�;w���r��uYt���tW��( ����#�$$Br��k�2i�wY��˾�/8����Q�f���U�K@�=�q�U+�旄��y� ���!�E;+I�R��<�0��������#�)p(��R�8�;�*Z�h������K�U����:'�������NL�0w�lc�Y��{p�~ew�����aL���di\6��T[�￴�)��)+�M�S;l��Ԙ�tSI���/)AN�G�2�j�
:������Uխ}��m����}�Ԍ4�m^^���-	>�u�`9�1�TTU	�c.�
Z��tGo	D��Z�a�]*�?����
���ꪾ`� �ǂ�y6V"�]�DZ	���cA��Ħ5�?����H*�ebJn�a��Tfe6b�s���UOq4E�0��+?{r7��ER]���J�́�΀�?z8�]%�����}�1G�*ZA�$�b��ho�}�1�uNc��ٌ8���u�g
��{��"����c䠢m�-��+Y>��ꁝ2���$���f��G =� �
�8ŏ؁8����=���U,�����j��j�a��)�>��ʈ&>��0�:��撞Y���Y������F\�sW3{+�&O?�I�P1dD��0Ǵ�7�C�Y�Q�o��g�
�>nN�'9���LKn2��fk���}6ҧ��^%q�c���jN����*wM�aDSΨܚ��!�2��vQ�B���-%�]��N�P��]�s���ZB��AY���Q�2�}ئ�D�icG���i���wP%/�@�Y.T�eQ����#��\z��Z��V������K�(� #�s�#�@�!Vz��ﭭq�Ȃ���>
� :�L�L���,~�XP'J}����_�sSV�'�P�O�L�d���W�t�z���fB-_���'r���f$�����:'g	�L�0_��5~�oO��ǋ�E�J
�"��=S�50NV��b�z{� ��a����(�T��)�=�.�Q� �e�%s	���h���I���"��rS{����X�)D����Ѵ�28���S'ɣv(�N�C}����c�0��K��4[NO��g�;�0��j�ӈT
��b1��i�Y+���p�i����ۺ��<#`�O�6)(U�ܔ�a%bO�09�s$��)��ܬ��*s�-�Iv�ҀE>�C&���DcA/��y�a�$UG�Pz@�.���29���)6^�v^�9 @=�V�����۽����G�����&�E]�A����]�`�N���`,C��/
�y�L��4�y���ꭲn��Ml���u�5vZ8�*گ뚨�Yau?Y'r�Ŗ��r�"��3��5���=׌}��b��#q�xT*8�nAOmF� ��7ف�c��C��E���ܿ�p��a��S(���ГCd�W��L�]���E�/�hcP�Fò��)����봅*�K?;k�Y0��!��N�^��恻���<&+������y�%0���/����Uk�������A�OuX����=^�9&����?� �r3��U�6Oו<�A �]�g��(vxqO;��M��v� ���B6�v��BVl15w�ݣ0V��`���,�?��2ZA)�y�C�2��eT{��7T��bБ�ٽfRN�\Ji|��0z@�\L@7Z�7A�����d��1�:¸���W�Ý�p��e��ei�B+M�;a�>�9�BY[<"\�9��[$�2�/�3Cq]��t3�ߗo[eh����g����	��n�S ��-�0xɁݬ�8<JE�)����&����L?Ow�+�t"�}���Ƶ}=�*����WrWz��3�
!�)С�1��8B��9���$7ɖ9��1:��b����k ����lh�n4n1���Ux�џ������f��j{��KBS���YU�w��l"Fꇪ��KwV��ΈL`ƙ�6K$�|9GR�6���U.1nZ���)����!,y����[:�{��"=��w���/#���l�V��~�Mau��M��A�Y{�l��c&���C*IM�r�Wn�E\���-d�}�����C�Hk��T	��E�8�=�=?h P�6	ϊl�NhJ#Gߎ��	�繦�+��D����s�WPp�7�K��T����)�*�ݮ�Y)�a[4�����1>�_͊�q�X)
�U�!s�r$�u����i!�AG��Ц���A2t��Үu�Jݒ���[��t?��&�<s�;�wd�P��I��G�
`���Gm�E l�1�	���]Q����$���>�SKʍVόP��Hz�ɰEՠ"x���ᕭ��s�*��G�R��A�^�#tb�����S|g���_��.!�AK�� t�{$�7����>��Z"�W�.CS'������� �?-���\RI6�/;���;�>J� ������P�1��@` �n���$1�?����]p� ]ϖ@/]N�X �c�8�2ć����,��N���=4��>��ES�V��&����5�ArMO�`���ZD"0]6C�zcm��P���Q��Қ�E�0�ڤ��x��gx��'�)ü����&O��ja�^h���Ϧ�6R�p�vs0�s;����R���v_�&KhO�|+��wHl�i�=�P�����*A({e:b��^������B���qC�,|�-�~]�� 6�a�^�!������-~��[��7�i�B�\g��B�*��uW�C݆v�*�T�U���-�;c�6+��}D�a��ݫ� �5]�!�vm)e|/U��
+o7�� �ޒw���M���d�cf���~���L��H���@��U5��Ѭ��/-D���_�p��lWfZ�N9\���:E��m[����ug:i������@ѣt�p�S�
�Tɧ��'�I"�yvue2~�9{L��ϥd	J��� ��E`Ⱦ�p�qHH��� �)5`J� �UdMKk�c[ʣ�&ݖKƞ�M�j�\خv�*�mdJPE"%wTY�|^U�������Z!����U1"�cUw���c�M`�zl�l)�{�h��"p6(���m�8Wķ� +螀�}+F������&	���F�5B��c	��'f�����.3&^C�X�g�7M��M5tA��$I�ZB�ǐ�O����m��6��,�hH���L�j�ST�w�D��-rJ2�I�(������jj3��`��J�ܿ���Ğ?�!�[�M����V�iϧ��t\i�BK<I��[���7!�	�d���ɒv���	)���A�J�}1np�L��Q0 حϯJ�|z ތI�o8���ip��w՚�_��pW���b�&Rﻳ��'�;M7.{�2]�Ï��$�M�*wxe�M�׏�Y�'�����51��$��7�|��P�rd]
�['k#���N�����	%g�;����ZQ�c�?�*|����X:~�q��,�y��geU�5�~Wy��m��¦�;��ۺI"��Żw�c�g �2"�R_��ӣ-�g���]� ���:tΧ	E���A�?��{�8���{Ľ�r����\L�!������%Y.0���]G�6��6�M"������[`+t�o���FV7π�F���~�m}r:γ��d�y!f/�`x1��w �jC>�܊"
q�:O��Q���i%C����<��*�GF� b���wطlo�]�A]K���2�vb�P���G�_���
��B���	w�Kp�+���%��P�����=+�,�vo�V�O���mk>��&�dmPS#*Hd��wz1�Sdx2���O���Q�/�dǥ2�� ���۸o��NktP���`�č�f�#���X�F��7ڽd!׹u���䘜�%�pw��MА]h!�Pƙ��7g����h��p�B%v5���+o븩�?��+㑒}�^�����=��DsTМ$�U7�ǩ>��S��)�̠�,g
9j���ڪ�G���Z1���yټ��R8Թ$?������P/h�"d
���Έ�`Z�W�q0�Wq��=G_ǐ<od�8�{z�2^¡����&���I�6S�	���mbR���Elb������u�206�.������?�3L'� w�7N�A?�U*�J�˹x2!3�i�&�?�^V�@}ݓ��a9O��Ga	�]5��Tgt�kd�%�X�4;�!���𑨖�r���}W�4<Ŧy�8��L=u�����	�A�w�8yÐ@����L� Sԅ1֡;��>����Ol�)=�x�9�~���߿��5�EX����aw�[�H��R��&����^�_ �{s���`b���{gk���G8��2��5`M2��;��QSN�;� ���/���fc�P���P�b�ӻ2�x���rm���������l������:'����z�#�rdqK�*��V���kWa�<��JoM5��IW���G&A�$~ʕģfg�_}�창��;E�"-�Nf��<:_�s�+f�/K�j	� ���M���hO��Lw��L����1�E���}Re��C?�m�W�@.���'F]��%M65�~8E�{�D���j���5<"qw���>�`�H�$ 	��9H�dfc����{[��Wy�Y�p~�!T��x�4�F�a��rL[�WRѥ`���[�;d�	�OqJh��#�w��^#�ai,��ˆ���Z��\�xt��u���j��!�2I����s ��2����@c^��+�������}����S������f�{�X��2ĥ������S��T�%C�o�esBh y���F��R�$Pj��MK�١Wq��[r�EzX`/%_a�	�n��In�<mk�A,���ڎ�0ݙl%��g#�'B�{=8�Q/���[�e���c 3��������J�P�&�pv�g���Y�K(����v0u�K�C82v���ۑ���i�ՙ!q��ϫaZ@�.�L6M�R��J�im��?�U�9"����rw%�vW�s7�[�y��y�!����?30a;3���'�\�Xi�п7�L�IB?��}��E���c��&-'��ee7ٺ�/��Ax�8?��j�����/4!�
Bs��� k��`�0n�4/���(*B�uE�i&�z�p!��'�-d[�&d�f�g�"�VA�eYU��M��}��n���ϒҵ�#t�M�?V;����cws�԰e���ʓ���]�	�!����uH�0�l�5�0	�AZ�P7��p����r;v��y�H�G�/uU��L�Ja���&;/�?���dԣ��F;Z��O8j+z�¯��Z@cqz�v���+�r������v��ۋ;~�w��n5�|)�{1�6���{�vth#�t��iN���b��U�=���G� ���vaH�7�$��5���iS8��z-�!�]��OM�^a��u��K�����������澸26�]D>���B�_�w��Yc�F�If˳��1��:O?��[X�o�J��zH�K<B��Zw;�\t��}�u�(�f�rH姈윧����g28�Bvi۵�\�j�P����$~�w��P*�b�@ҿ�E,>Kg���'���@[�DؤԤ��G���U�#�ˋ1N��;;��fiɓŞ�%�8r���0�e��WUi6
�Xg�#^1���^ψ��"���f��(��sPD١ŖF�ݱR��B��k�;�	�&���*IH�����L���\��w>�@=iBY�Xm�<��;��4�,	:�cɻX3�O��1���q����&�m[S��|�χ�_dP@m��K�C�rnT����o��3CN��Z��K-���y�� r]�$/^���,]���(��k �*˶ &_�M�ݰ���Ȑ��l�K�z,�+)d�&�n�Խe��|>��ZY��[�|�/Ȉ�6���(����l�n��3q.1B�� ��R�TQgB�M*���#�U4v���lq�I�ٌW'��v"�a�Ѽ�����<?���$"6I�Ux��s��J���2FЙx�c�f/�Zq�1l���R�Q�Rn0i��9�:��7�{��=	�Ԇ�u|TMᫀ�����X�Զ���0NeS�#i�O����e�u��Z���AE��� �ZaႨ ��>"��I�*w<됖g>�*��x�����W�3����w���qHd�p&���O�Jh�͏-�!kTk��	m���ۄ�楕@�r@�!��ӁL׾�"H
@w�O�}�B��tTG�;���|�ɠݭ�*nW��n�2�ɠ��|�@!����k|C�%���jԖ��Ļ�d���Q^]P��H���,��YuM���1�?k�z�ʇ�؏A��W�K7[������:�E�:�bFH�#Q���+QtŷaO,�����eÈ̄	�Y:��<�%s�FIf���N�W�$ ȥ�2��-CV��p8z����C&9��3Rq@0�m��Xy7G�^�c�Sp�f|��B:Ī;X�e���@o�P���ڸ�3�c��r�����;��!��Jfa��׳��L�"���u��#�\Ty��J�We��:���2�u��q3�L5����Ah�����:!���3�Z>��^^k�`���oq߅Ր��T1����*PS�%�bm�� e���)�}Xu��H�N���#L��xf^B�O`TE:���/��(��;N�Bc_B\H�9r�^k�S��=�጗��~����IM���/���1���5����ߥ4�<���#�%������G���O=u��t�HYp��>�ufgy_�������)�BW}I�-k�7�/�.�� �r��5T�\-�F�>o�憴m��5=�yaZ+ܾ�a�4�8���ߚ���I.{Qp'��Hi�6�Tk�R��K�dZ4���A�M�0��X�:@�����QP��k+�yU�+)���fI���ŉ��ť�C�E��������N~�-�fE/�����m�M��؟����]�)�������F����o��~��\�p�t��U�>�P|ߚl,�X\!�g�=���!����}���$����	"���
��v/�]͍}���o,1�A�@���R� )[*�d$�U)�P0��ETu.��e�	B�<OO��i2�ʡ��f
��G�M]��rE��*�����&�q \���G���&���K�8Tf�(����t,5�����+��$�V��n�y��]Ao/�19��j��Y	�Z�n'񥆏�P{�/�9�eh_r{�Ty`���A����Fq1���9��9�P9��g�%��K(dt�vez��*�~�/D:k���+ TyP�&�MKީ9c��eY]��h�۠��^E�肅%OjU��m2�����3�U�����7�PmAM����}�	���,�6�7�
�$~T����`�t�h�(�o�p�<�����'5{G*»t8��~�a������b�I_7�!�acS)]u�,���Ӻ�X��щ�&��l\Sw�2B�G,�f~'*b�ێ�`�y�6�8�%*ˢ���|]:R�O�	$n�m儞����� 4x��\>��q��I�뚥J+�,����<UzƼn�� �� 7ѡ��y�Z#7������~��{mnЬ����M�_:W`l�w�����u�t�"���Q2���� ��[ U��7�7��(EƇ~�����,�b��`�_t��'�h��}�Gؔ�<�����".����%g���q9|���S<��� ���㈱i�x�i�_q�G.D
BHu�����sTaR4��s���+]� ]Q�iz��W��~����OQ+T�*vCf���ɦ<q��@��L�>�d;�%�(���	� Is������tM��ٟV _Z�ũ��3\�j�I�HtK8�H��L�'nk>��p��a��/kQ�������������4��5������f��n�P%�$<����\luCh��VS��R��&��\f��K��~+�lD[X�W��0�H�U@(׬����}E8D��iFv�25�p��'>nut}%B�/�!o�]<���f*l�?i�L�B<�n�Nˤ�E+�����m).��ތ����9"##�|��A��+E����N�y��?Y��^(|O��9�����!��:�qhv���l�7[��D��w������P_���H��y�D�D�u�T����5�Tĝg]t��Jc�TܤPЎՙ
`��u���6���nwݞ�dB����e�p7U&���o��<n	W�T�LGì���`\�,��R�gP�Z�O��H˰�'�.��pG� tO�"INu9|## D������	�brkѩ�	�C�m7��L۪� ���|涚/��	7��is��?i��������؈�����m�Dґ��n�~A�WN�Y������\h|G����6��Υ�-���d��m�E�v%�*�N�$��ЛvC�R�y&�C��p� �`VX'	�l����U��b��'
�=z����+��HƳM�ŗ�Y���F#�BHVQ��u��\�Ø���"E�|:]2���bئ����q܂ݙ>{���1�\c+-u26! W��0��E���h���g##R�r,��b�_R�y���U�}z�V\Q]j�dm;�N��2���s���N˔2�Lk�_��yM�Kg`9]��s5{r8�\'�$�/�Y6�_ݽW�?�s"��Q�y�`�0�7�Z��:d�fz~)Xqq��J~&޳g�0�]4�y�O�9�3��hr�4�#�ϝuY#��X�t&QJ�G<%s�8����%�gq�HVbd���R�����7Q�@������m	�����{��3.4���}ԣ0�? S�sK+|���: �	� �Fc�bQAY�ͼ�	��۔��ao_�����+H��M%��$�/`pЍ@��Cű@>`�(%�!Q���$�������������� w٘�r�/C�`��!�75�}���L�Kv�4�������$՘�ᬏ�W�h�N���klb;�=�/#m=kG�;?貫KO`�D�E*����������m��a�+���4��4����p���z�`T1���r�!7La8�n����, `3���'�%���9Q��I���wt*ѕ6�������pFקE^JN&/���K�~yj>L�n���Bc�x��^��"�M��>3|F< 1��\������	㠿l�dӜH�ҬB�.��wh�I�1���5�ex�}I�8lj�����q�vxRN�~{�v�g\p����U!u9���m" ���u�w��S�:��s��k�qH��b�Bm��!�h� �ś�*tC2nPh�4�WPh$f��|E�9~E�I��5�5�"R��ū��X���;�:��@��I�;S߉oZ�3m|/�Le�����? g
��.��Tz����viU��{Ѳ0�}0�/��tR_�]�z�K��'l�]�d�"��p�� ����>�@�u(�ཿ��$.�m
�`\^���鹖��|��Hψ�R�[�[Ft���uY�3"vϖ���an���K�{�]~�Φ�#.��I-��Q��W&m�a`���,d�u�)P�Y��۰�u�;���(Bكh�vG��}�`a��9�P+���R:��6���?��X�	9K�lq	m�i����xok�J���ӱ`ģ٦��.�~U��(R"�N� �l�c��������*��p�oz����u�Li+�ƩG�������T\I���[3���"d��3m���v����aQ^p��u��iH���}��r唸BiSg���9I�U;F���N��&����fG��j/D_�R��G]b �GW�X��Q������m�-����7���hz��GK$4��R���o�G����w|[kzf1*%M΢]O����~��ӂ7]�?�2��b��s�@6�U�\~�۾��s=�l�i�A��j�5�Q$�Iy�^tGs]����y��|�����AmW��L�<�*D\�W�׽EH�x�3��������+�O�S���+i+��9�~5����nˌ2�WO���e�׌h�x�!�4��B���Xq �Ͽ��|Z���Z@ I3�'�.@�	\$!�=Q%�hH$zY��}��F��#�{�X�r���f}(6I�(�z�-F3 jZ��_v�4�kOøG3���q;(�v�*$��х�����X�}�b��&�8쏮y��܁!��l��3�-�Z�$�~ژ/FG�C����L�*eX��@/�&c7����R��d1x��I�������L����W�J��v�Zdz�KT��Ȝd��3�����/f2�5�q�.6�R�!��SrXc)lH/�m�]�qc�x$�2>G �|�e�u"�s㬐<34�뒴��̇�݄Ǧ���l �O�G1�N�c�q�g�ؽ�Y�:V
D�rF$̼����` _�8O�TL����dE��Zj�. &"<ZH��1�� �-�`�-���<���R7��J'��6�f��Hn{d�DC�[]���D�8���{e��:���
 1������R7̷��O�e ��H ��F������̀lkp�׽��|�}s����f�v+�3�p��r��[�����^v"��]�u)a��z&T0�J�E/����}�&8����s��^�c�N㴇�An�~� V��n�;�o���kJJ��)�u��l� ��i��~6�&�=$����V���E�%!Z2/@b��bX��tO���$['��UŁ̼c�p�a9�W��h�b�pfb���V'8�͹tgK��=�@P::�32Qv�4������d��o�t+�G�xH�Q �Oa.�P��Nq�V�KVY�2�>�z��$�3V��ŋ� ��lR�&]��G��l���|��M{�
�7埿�ॵ�mmr�ӿ��wY�#8CG�%t��oi��Uܿ�2�Z��li���樛�_$��sv�2{�l8��C��^���p���$(�?_7�>,	>�����L���/r���$�f�g��$	��}O`�3'N�`8����f�j�Ro�8��y���#����ݔE�Pʬ�,JS5����ҝ\�j`Q�9m֩�ߛ�\���[�WI�@��_�H���wVu�m�!n��r\+I*yСI��g~�K>��<�B���Kk��@7��������}x�Wꉈ%%ѝ���k������2fq���]I��;sR-XE>[n�8�$Fl���M�&��Uώb�ޟ�>��Y�C^/X���vC���ͅ*���U�������AܧKTE��g�L��_6R�k�ʖ{���V����3삉��_;�Y�w�b#�7Z���ǽqہ~��(��&���M1w��*�tݓw͔�;n�5�
Ϸ��p�gF���6�3�	t;��W­��OyQ���H�� �w_�j�i+݆�TQ������P0:j5D�#�dzv;Y$$Q�����;R����b�i�S����'V���)�+,)+̎.�Z>2�J�	����2�� ��g��iV�������u�Ū��ժF�R¨���o� �դ9���[�g�=l� �JK��E�[mۚ�馦N ��5�k��+P����cA����}k���K�c��Ã@��1����Af1S5�)�����
j��!3�ȍ���_ӹݨ�M֓�؜Zƅ
,��{��/�΀�X�aO�N_ϰ�JM�~�Ơů�]�=���p�5P��ߌ)^��Y�;[��6����(Oˎ<ch+3>���m$�* Vo]NqQ�c��I��J�����&��Ye�^-]S�Ր�=����q���Mz�u��{�_�N{��o��q`{_�w���V7�������MI9O��A��L��.k��q���S拑�X����e�hX�Ԓ�t��Sq,�F�^�����4܉�s������z'�p��P��ĵ����J��+�݅8T��w�=��m� �oT��vp_Xd)��?����-#4cŹ
�uC|ʡY6F@���]()�7���\�<�� �c�w������g���\�C�q���µp�Q�����O�9Ȼ��B�����hc(1�= !x{g9(����,���w�4��%\��%�1|G����x�zUתx!.��]����k���Mnū���g��i(N��/��WY��w�4�d���m0ܝ|�#<�uQ�]�����0*=�����e�CF�-��ӗ:�(Z��8�bk�����:e0�������s��z���J2x�Mɍ��8ļ�r�Q���۽)��A���[�R\S�,X��(Z�4���:u^*h,L��1S�� j�^��֘���;��%nD���e�q�ؐ31�����r�v_�~��9���oG��U���VY�QZ.T�
Q�յ�.ƂlqC���6�V� �Ġ��)J4z�66]�V6�[�g6�^%��~���Smx"4��]e�&a��iN�Rh}������Mq�+�2�7�Z'}�&sl�U�,~��^�Gd�v��dE{�"w9�e����O46�|�	�Sw��Ζ)c�v \d��p�g~���i�*�΢�@�ܶ���Zg����:¿U������G�����aveBs%�H1H����X���"�=0��r��W�$]T���Ɵi
�t�@(���'>Lg��=��}�R��8��Y� ��p�]��>�R7:%R"�RG㴸i�m1Ӏo�������ѩ}���N�RQ�=��G>��P@&d���̇΃u���$&�	i�Ga���x��Wt�?��@���+�b���N���+��G�S)�%Fe�%��jn)8�m�o9�H�����#����	�(���^d؉4{~�POzi=i�

����]2�'��|�ڪx�L�"��r��5IL�G�n{�~)���z>�ц�'?�����qJH|�E��Y���v�ϫ^R�+/���J~�V! "Ӈ�5���_��R�c�̚X���լ5ʽ;���m����}\Y���2Ϛ!F@����� �6XGZn��zfk�t�2����}�{�@�Z�6�>D�l��=C@:�Ik�b�_�����D��]���vj*qќc]�[�S�W�U
����Z��#�û�U2ra��G箠��(E�5������N�j�U��MT`�W��隃���żym�K<<��'p� �������y�w��n/w�%f#B�3I��5S��O��{�e�P��zܮ�f��L������-��T�0��2N^G7*���}%�;�2�
��8�G|��wV��%v3Ztr�iիE��C�7!L�?'�l�%#2y	����8@GBi����AyV��d���N��-�A9T���/�4��M<���Z;Z�����ul�'�*��}
o����A[�釼��`&�Gτ:�+��X4T��ZD�&�%32!��FkN�8{�(�dٙ�/w�п\�I��`J?�h�'W��$�ܬ���ĭ�!�m�P�x��t@-	�!PgՍ/'�g[��((S���ymj&�3�3��=�NAE&,��mu�} �7��@36����}|K*��S���'�a�F��L�eA�$?��2Ӿ��c�m��x�hjT6H�]X
�b�Ү��9+ qe���F�����yz��4����$l�L�}��]5��~F��y���ީ�myQHEĄ�N��~�Xi���+��W��2a��!��p�&�<i�����	?�~�QY�W2�L�˟q�*+�<LWi˺�����!�X�\��O"���Hy,o�}��|W�Z/��g.��DW�A�i˅]�T;t�--�Ȅ	I?���m�c�b�
<X�f�Nk`a(z�ͻ�!���/�s7?.i����`���&PB}�`�T�N��������!��d݆�X־1kT����b���\�虍jЩ���g�4���%�J�9UbF�g����8�E(lc���@6���q����5[��Z.9�=�x�N����Hj-�6�`2�ְ��t�I��1�vZN�J;nÇ϶��J	\j |Ĺ�Q�C���mWu^ ���&�����������%�"\Q��Aw3�	�P�ˇ&�&Sº���yA�&'��C��Q�)L����a��[�a'�����GB��]��,�BD�'�S3�=V�Ǳ!.ѓ��E���'ɿ]*��&P�,�W�"/����M|u՛��e�^$���k��*��_;�	�j�C�d�cX/���\�#2e�eRI��"�Wp�"�g���1t	��=ǂT�C���1�������ZN���˰�:]N�d��v9+x.r�`��#m�T&v���*�����NF�nϔ��B�~T���E޾.���o�Bw���}��~��G웬��.٬O"m���lF�*/��
�#�I.��`�H�HC��C��U��uaܗ�t�ꉹ��{��I�~c�4�2f+8}ٴ��P�KN��"۾0|D����3Wb����<X	�����_���~��{�9���#��ڛ}
�qc���Ӟ�o%���EB.S=��Py����\sk�Y]�vhT�Mn�T�Eոt����xT���O��#����X �&����v�ʐE�� Ҹ��g
�N.�ԥ)�7,N���5�z���O/s�U�nņ�ߏQ$�za� �� #~��ȧ�{��V��.b(�����Av'�^�զ��ߞ�fe�>��p�1]	aJ��@'x`�oظ
� kV���y�k���k��-q����nu�D����a�R,	[�4����!)֡N1?9��w)�U������p}���g����]JY/�y��|���7���RS��<��CK��6�عحqg�Q9�ک*���z�:\sϨG�)u2�ε��X���^�o鹽U]|PS�KǄN�!�ƚ��D��i�_�I��\���ω�3V��g���뉫���YC��6��a7T%��C��
��su�zќ��Pm�{�sq�K�9��M��e�� �E�>δ&�u8~��fX��K�~�Ɇ��\.C�cxM�h�mF�
[�Ҟ�5�G�=ϒd�Z�bo��� :">�t�~Q�FK		��9P�&�9zO3���aa���W:2�]�n&Cc��PK�E�	�Zp�
J,/d >�+h'5�(Z��*�R���gJ2t0�∥5��)��i��#7[�ө�D�l?���6	{�(�)��	\����\0�����d��[������d�������bKQ����ti˖�s�H`V�M-�κ�M�D��i��3���Yf8t�|�|&����^!�Y8�L72%y4�{�G%��%8�
�� ��
�I���3�΂$�Qʣ�R؊C��xߣu�*��鉛7M���B[�j9P��8LB�y3"H�(p�� ~GB����дT��:�et�6iɹSXì=:�����]�LA��=�~�`��v0�w�pw�=;Щr�N{?X�b�l�P`����1h��Le�(j��
�'}6�<��J7�<�7N�4�<�V�k$p?�I�CG?�]�����G襣Rl�H2�]��;�7k��Q��놎�qp�8ߎ��>�u
7F<���E�9,�
�oGLuKs��e�< �P��a���Q�/Pwl�@��^W���,�U��~&*Ie�d7��R;��TFn�wÕ��"s�E*���HZ�m�!�ݛ����E��=��ep��YX�mԷ������f�PnNd(W�f`0��}��R�T��q1J­ �/�/�0Q�"�>ī>̆�x_h�x�<���f�u�+g��t�v�����	FnK�.�mA��$ET ��b�#��U>"�LU�R���ͳ���$ΗLV_[I�SVU��>��"U��c.��M؄ǿ� cL5�;ᒆ҃ɊR�������<p ����0BA������m?�j��3�:��6�-�y�ؕ<��"*,�ѺӇ�M�)���Å)Ҟ@z.
QP�;C����8�S�`�9L�|s��0�̪� �����E��|5�`t����v��!������%��0��%�)�' >�����M�����ky3�ԸR�"��c��o��`�E�}��2`+Z��`'����h��5�w�T�4��j�-��If\��Y��nci�o�2y-�xz�TO��Ժ��-���`���T{�
ƺ\�����??��H���A�?�eڽ�ݣT3��L��P�������&�*�H-.�C��H���mK��û�_Y3�$���lF]�\Z����{�˄�!j>;��R6��;���z�B���^��,��?�%�	uI�W�`/S���RM$��pM��B ��H��kIx��kV�%�g�(E?79�eV�~�MN���7O����DsTi�[�p��h�N���n"!���$�3�����Z��=��1�V�%�%���|�Q{��o%yx�x��\X��{6n�ߗ�ݗ�����'P������({��Po���z����Ъ�kj��R��|:�I}I�h:
��>­��$������
�
'm�n�&��#�ur[��X5�Q��!��R��4����hV���)��6Z���&/��D&d^�Nh���8�Ҁt���r.+,�/BO�GJ���G�����sY�Q�;0b\v�h��HC�8(_��F�U�#��֊���?0ͨ�����'g��q	��_u����=A�)����#T �;7B���Շj�� mԳ���L����q�;f�B�w}�y]`Sժ)���!�S�(��T3�����2xϔ�0~�_���#���F�qm�V[�A�_��>E?�����&�����"Fc/J$�6øݯ�������l,6��am�y1�t������[��P6/��e�j�̅�_�h�U��T ��]�g��t�"	?����f@V���i%����,.��t�7�����[�xٛ���Ke3)T�h��3.�R����R��I�f�η�f�@@�]̀.ӛ�X��?!�o|�����:�{�� &�
,����q�o�w�a*ɩ&$һ����`e��M�hm��/����1ذ�C|���l���0��k��L~[re�X>���q>Jㆋ_R�~��O�;�99�|�1CrG�d�1��?�3���J�խ��9�(ñ��� �+���({��7x�^X�G"&��`��s���1a��bB�)�\�<g�X����D�jV� � L�T�F�������O���;�\�G@��Af������V�1��]J<�J�C齩��I_�;�љ/tG(HY�Cƹ?ĭl�C����AU!���Q���8<���ݖ�+�Sc̫&3�H����F�Ph�@Ӗ�%�j��r����Uiܜk��]��,�X��*��7L��uTH�|�M]�&�m�_���^ɶ\l�Uq;�R���-��!�Ӛ�Bx��Prs���o&��^)c����͊g1 �����Yg��	������nՍ�����`�ze�e�+.��,�1,�Z��h��ׁq_7�rR�y4i�ѥ���8���S9l,��"$N��&E s���#
Ҙ^��*�(�^�%�m��~�,��DU���(񵻒&F������i���}��\�coC�����:*K���C����nM���j!R�� ��_�,2t��P��7�����1���jM�&�u�bc��NY���9F�S���2We�mW������eO`��ė��#e�C��
)r3Җ>�;���Ei�t��&��Dj��S���i�� #�~�px/���t��v�v~�e$gs:&�H�D����.�*��c�sP0����P��g 7F&"��V�d��X�M�8Gřk��4�FM� u�l�����i�"�P�VXO��w�.Sb��aiҘ����S����[��~��~��goW����w�x�]��l�X�2�2T*t�`�����hT�+�ZY��z�����J��K��erF[&��B��N��!�~�1q)�|�B��8 x��o:����ع�dC�Hu#���[�5�z[T? {�g@�
5j��#,kԑ����2�Sٹ���q�����Q,�'�w��2u��i?��
1d�N�>"�Q��q9*��R�J_S[��E$a~��@p�0�HZ�rz���1�~-ϯCy��b���~�SS�t���g�I�7O���"��x��B4��YQ#�gr����F�_��R��w�|����I�}�j`=���k�za����V���z޻P�/���2����S��%�|]"F��n��6�.�=g��ZxP6Q��x��#{ZJU�K|%|��Qǃ�=�m�O�3ݹͮ�E Z����˕d��Н��Јg�O�1j�Y���
��~uК�CF�������
G\��z�HC�d��*\�b���M��6X���F����������)�m�����z�h��/I����Cs�ᣰ\*�Ħ7SfG�ȹ1Ԡ��u��������//���ǐ��{��m�(����X���s':̳�����t�1��.V�Bؠ.5)<�������=IF�Ro7�Z��׏�@�.lz�w���A��`U$�B����K�5��iɜ8���$��A[��9)m��{o���Ԛ�iIW�&&`9#�v��Цw}@�UO�ڨ˕W�G~�p�T�48Z~EL���&��k��ԷΊ?n"��&Є�wώS/S��N�L}|����	����� (�5Ǣ�'�}�����/�`Ҧ�B򕠕!���JU5��B���]�>�@��}��,=��خ������潏���7O��aW��.�΀��,�p8@��m5�&����i��j�d���,E�u�\١O�m�1�`�0'>�4:��k��M�?�ж���:6)@���(����^% !�)N���Lc�,��|��53�%�+��v-�e��~y�^Er�W#y��ꮲ(��[�Ҍ8��;��Y��Y�v ���P�j�).�W!�g�)�!A00K����Mαs�o�
�z(QO�՗%j�6HD���B|g�ywdD3��r�"��������>5� Y,�=d
I\1����Aq��;8{��1��u7�z���I]�FYUH�����(j1;bd�o�mzǷt���⢂t�?��f�M���r\8#R	&vRe(.+B��9J������:(n7��e�_18�<�w5�?��HO�K������F����lu}�i�z�C��>���w!�����`#9�������O��Lp@��f�F;'�2�$y�����Io���Q��T����j	����=?�0u^+*=��\�'z��Xe��Vs\�Tf���S�FV���>ݷ��[
	G��1QoB��l��.���3��8g�ȶb�ŗU\$��p��κ;=�!��U)�D�X~%����w�k�����<�{Ay�kH^c��f��1h�r),��V��@>��pO�s�n�>o��I�k�ىs��o���me��"չ�/�{�D�R�ŀq�+n�2>s�?�(m5
��PHY4P A�֒�`�el(�JZ-�c��v��Q�;-�0�|� ��$�w��($�%�};B���3S��������`<�k��r�����ޭ�z3�0��������,�L�����4����J~ȣ�4rP��qB�K��/�}�}�<�>��V�Q��� e�����\"I��x��rdw7"4�(H�0�!�Pn�>���� NQ��[�=f��eh9d���>����� g$V��aN�$�MFb��GH�_z�j�θw�4��mg�S���$d^�.Yd�_�~O�/07��_�&���i���.�#!1���?U7�J����p�ݹ0�5��-�n���131��݆� �։]��v	��x�^��K�d_��|��ޜ�'	��-��=H��³xR%P��������`.�����|Z�G��(Ӧ�Pн����z5.�0N
Y�9����[�#`�֠2|�����۩'�;�@Bd$*EW�/�s�/w���v��%�x`�@� Dz��_�
7��L�䆲�~Yt��L��gi�e�]�R���l�&]�۩<d�s�k�#gK-�"ml��O����	��+�y��<��7�O�´��f�����55A�n��ӽ��`KڰD 9��e���E{&��%gu�9����^HԸhy���3b�>�_Ta����\x�iO#�0.�������`�.}Qp�;'=�Y|��]ouz��[�&P�����kL`щ�@S�9=��9��a��]v���~䑁h Pr����P
[�ڳB ��q���j$aұ�S�ح�=7:A�Y*s$���1�m$��(�ޮD��ȗ2��q�:|�.�e/�.�뻼���X��AjM�W��ǹ�P���bMxGq*��v��;�Q��E�|��Z9�ȅq�f�VkZP���>���+�tZ,��k4�Sdf�
��|�)/GF��}Mߒ�
�wz��A�n�I1��V,�B���3��u	������f���W� $��4RL�sR�_<" �7���B'o����b�x�J#�YU�6��p.Cl���3���eQmΥ��ɭ��nu�1�E0�[|y�+0T�Y�I�ϫ{��3�۱I�_~��~�LÒ�����I`$쥞֬���iJ�y`��03��
��ͮ��`h�M���E������� �Qϩ��iC.*B�E�$Q��	���_�@" ��t��c]��P�M��d*4Ds����\,ϣK��<��>�y�Ii$�HG�a�e������~u�������B�~9}u�/�--�6��9�)�a���~�F;�l􋡄f�4:*�{�6b�sϫ������X�°�B�����a�݇�����Ѧ�2�eu�˻-���e�DPz��6h��t�=vf�]�e~�����zฯ[=3��	�Itǳa���ܽ<F�V�Q���lXz��K��_�f�����8�R���bj��a 3 `�4�I)�������A�1aN"C/�Vt'E��D z�^o�����xhj��O8d|�J��Z�͒����^�R��d_è�(~zԷ����,�,�s�Bk3��K��$�ݩ-*�g5�S�()*n�ؿa+̰���.���1�_}���5��Ӈn��k?��9/dk���Mf�a�T�,i��kk�*���4����r.;������Q�-%�Z��:��D֬LO��o�b����%�?S�es���~x�铸t��7?��B<�3��=z0�[��.x�Ē��+xI�x�7O�B}�����U=@1�:Q
�$��h� w�H����6̨�BΝ�H�$�w�B����3�wz�X;�d�10Ds`}$v��2��Z��`7.�����:��9P�{�h�}�&�6 �D��Ę�DQ�/S��R�3;�ԏ3X%����EھT�g�����z~��PgS����U#\��5ְ�U��B2d��U���*��i�jc�~n�<���Q;�*�Qd��8u@��|7 R�K`�p<�#�4�;��Ee/z����X�D����W�E�XD���D�fv� �RD�X�KwKp��u (�A�c��\z�?xH��A2��J�('���Q��O��<�$ �4�4�&����b���ǰ�юd��i���w�g|dy��7�ty���!��e�V���"��Tz��e2��p�L�����,�@�9�	!11���[�2���t~�X�NW˦���*�C�1K��:w�m��u0����Knyum,�CÔ=�Q�����:�54WP!oja= &��O���-������k�8�v?8:!��˛�<��
M���A.^g�Y����u'jZ���Hg��f�:@��1B|
!�B�ٞ�ծ-�2�xQ ��hq�	W���]��s���%�E�	�O�^C��G�6E�YE.5��9؛�������C~�.L�����RI3���4.<YѨ�O�[�`�*�d4pO�o�,��%����?�u�u���R=<b��7�?x��4�����pths��fEm��{�m�sA�L�QI\W�g�4��ėE���)W����F.�:�`����v�+�ٵ�������\m$ڨ����mP�Dc�//r����I���|�F���[��h�0�?U�����Dǟ�A�>��!`�}���Q���N��X��Ek�&�sf�L��7ՈZ>���;i�Vb�St~t��)�F�.�=�/��6�T��bC`�OI�!��8#m��UK���� �3b2��:�X��}i{{�'��X�ʻ�?Mk���9m�L�$�k�e2ה�s	bh�݈�A^ߒ�'|���R���X��Ξ(E�T`�N��'��'������*��Rt����:,8_���Qz���^
��z�^;a�d�¼��r��7�xK�\XxF�2��M���{��׻ �ۨ��f�~X8鑻��2���o����mp�2�G�?��6�-��2������B�ח$��2����5!$�(u,��H��iJim �y�_\Z\<8��_��E�r�[
��8�R��'�^��iGC��������w
�����,M
��ELMr�8Q�æ�^���#8�*"b��Kٞ	���Ο����<	�]���EE^� Ę�c��t˸�y2��'�����M�XM�ГcA:�������X����TA�Į�h7sh*���i���KOdq$�i*rͼ?K[���6+'Н�Z�y�z�'�س�*��_�s�m(�`�{G��0K�����avpBZ��BC��չ��_��m�����'�d|��I��FЊKP�6Q�N��~l�3���h/�y�H�<�ňo! l	�iI2�uU�x���G*�~�9q>|�����^�S0�\�`�0�
`�w�P�~X���Q"NPs@���K¯A�PU��N��jf�`>2t�!	��gH�``�Թ���~3�T7fa�ۈ�8
}�`�c|gk�<v����I�!�g��U���w��uRތ�0�A�o�hs���=����R5K�B�g��vZ;
��\9(�Bٚ���<2�^��v�<��
ߙ�9"��#�H�7����xX-T��9�m�q�h0�-�yʝ��X��(yu�>C[�T}&�7^5�D�Y�d�
��&��'�>Bs��+M:��Se���}{_x���h�P���ft���3�Q]�v�����_<��\�ϼ��҇	)�.41o���S��x{��\3��l�u-�H�HμYA!��b�`�q��1�6l��dK	UB��K�W1�B�CLk�mqb��
L�ƣh�t>��E�_�+~aǤ�(�v�$�v�X�.�l���[����ÔjJ�kϮ�! gCt�^7 $'1�T�]G��4��6��5q~Y:�sZ�O���˾�
ӍuH�̡��I�z�߿QI�i	Y�����ۀЍ<O�l9���. ���~�KUi��]��dc�#��g�燍e/v�����r�� ��
y����=A|1�j�j55����Ɯ]<��3͵���"��������帗�D�5l	e
�7�!��qy ����k�[1^���T�i�!��S�p�F�k���9ѣO�f��0eQI�+����sG�5���	�&����Hw|N���4�������G«3�L�:�|;)�z�g�0�9�p �0]A�s�5@��;����4� G���c�J�
s`�37�-tCl�(���8�u�WX��u����{NF����~�~w[��`�k6[Zsd�'�$k���q$IiV����0�A�G�w��w��K�P\6I����fP��C�%��ܽ9�xR22f�Ar�^!W���^B`&j%�}<<oM/��yd�9rKw��ˣ�1�/yS)���HQ@��s��f@@�+E��|�qpm�۪�97T�Jt9��U��Z��U:U�y�z��~/�ۊqXB�޿�bgHti��Eҍ����]kg�`�I����)������l��قeH��!�2��\_]#���ߡY�y�u�tj��ˠ�!+����p��5��p�G���Cnc��%`�D��>1� ��k˾N��H�O�|�= �}i�E������.i���-ۀ��7�@�3YuF'���_�U����覘��J�7X�蚠�CO�JW��0���2��f͓�Z����ZV՟�f�F㨄�� ��,*� ԸУG��1�&.�ʲZ�^V�~M\�\�Z�,ʩd�S���6�D������g�J��4}Eg�hO?݁I��Uc�?�Gv�$�b#q������=���À2Q��Ѭ�����Vg2�\U��U1C;�ϝ->�T������Vd�|6oq��'��������ǐ��z������5yIj�R�`W����.rrb】fmH~�O�Tɺ/
�M�-���J�N�-��Sjބ?�|6��0r��v���ӵ3b�C\�����Ń*��g
F�>�D�[C]4�}JX�
�;�%�C�N̠c%���(�:��s��I�y()�#�P~KW_F�N}��������9>�d��̾������=�A��zm��g?`���Dv���H��:eq��Q���1.�L����E��������R��E�S۵fg�L�?��Z�Do̟)���[i$��������t�S�4�K������M�c��קf�<�x�Oq �K&�{�CQ{j5B��e�S���}�n�l�dff��.y2�]��ř�y�}�3����tV���(ӂ���&ʑ䆧�ö�X���ם<��i�����!o�����笆�}�c*�Y�Vk
%=7�!s@��5�6쇽2|#��R�������n=~��H��c$��ԙ@"갹��^'*
~�J6���@"�R�C	��o#�wW�ɝP��F�D�?��ğ��v'�鬣LͿ�7����㺘�Hz���)n��x~s�@�2�Px �����HK��8���Tå:0Rb��9�g�)���I� #3m�y�PRJ�\7H��Z	k�o��\�g�G���j�=�_�6 �Z��~��)��R�\%��.է`���f9���՛�h�mB�F��~ke�%<�y�T"�<ʽY��Qy������Ј��*b�� <�3�*:q��~�����CZ�;>��o�*��}]6S���/�|�G_�m<Q�2X�5���~u�f�F�Ͻ4�V|�xZ�HHF�@.�f��kEQ�}��:��<�))�#b�ʯpqʏ���"�L��7�^�WV+�_8�~`HZ���+�6�9�gJs?�zo"1����P����R0|�"��ᄡ�KB(w�L�i���a<	���r�G�"�6��Nsĩ�(�Q%�Iy
l�L_� ,�b=�.	���>6��d��b=-��-��ĆZxU������aym�g,HIy�֦�?L��nFX�?�SG	\��n�&���MW~N$]�=++ :"�4���E=��xs"%E%�cr�ٻ'v����_��~�X#!G�|���'9M�W�����X3����6c��{0mL`w��{Ĭ��8�����!�3�� ��uˬ�ST�_f!��v��ވ�5�]#8hƦ������8��sP�ߤ�.�0���!���{�7F������VQ��j5�]L!��?{y/;�ek�υ	*��gh��m��ͭ�n,�͛�l� �~[��q�4}�}�&r|�^{uy�ց
�wV�i2_�����5�>�Fw�x�����i�x)���I<��+B'��� �J����s���߾L��")��\���B~�,�]�'�*{�[���V]��s�t�4!�9�d �	qc�\�����短�f��v�r�D�u�o�%I�52=��al�R�p���yE�$��|(FD0�:⒩��l��'%�v��@��"�W��dU7�֪T�,��تV�6?iKn�`�5��R���ѶzIb��*}�q����M��*g���%��X��q!�o��/���0��cL���}O�S,���|U��_�:}o��/�8%>���m6��f*�,�ܭ���
޾.�2����!��=�C��\�=�_��ܵ�N�x���x�c�;9	�$�p+��y���V!vm��X���V�pr��rL�4NB5��Z ����\AU���z��pfE=�����I�	��e�����^W_ٗ�A�bP�5��˶��1<�\���˿S��c��4��%�'�b�Ѣ��|��)\q#Ը�����(�#M��w��ӪW� Y-���I��4m#�C�?5g�.Xw����3�b6 ԋ>u$�[�P絗<�_mpkk�~21J��^��Q��B�ۿ�:Ȧ���	���1Ȏ���h8}��\���澰�Ӊ�bCa�+��_S���CھU.r�O�8�u�|J/�S�f��8�Ll�u�"�FS�6KQ.6�v+��!� �1�=D�Y�ӛk���F� �0d����ǲc�(' �n2j3��7����� 굄v/����K��>��_V����@�����@��:3���C��!�f��r�;���B�%���D�h�}�0TX!_[���&���2�N9�d��2��Y�]`����9�Æ��N���n|d	���|�P�L�������f2��͍���d1`�Ep�}qv������V\�(����069)�]�Kl�Q�p��$_AD�Y*4�-lŰ�Ǐ�y*��4{�AF������X���o(��"�(,N,��7<�����f�g�d�����[Ӧ��J��&�Mu)L7u柰,�@��I��2?�.ݱ�~�K����jq-�?��£T�P�Y[L�9)�p�����œ�)��ŨpZb��l[�	�K�S���b'�	���'t��0co4���Yc�lv�!J��>�E5a,��6�.t����[4y����5r4BN�h��ϨГ%��1U�5�AMWaLZ��nݨ�A-gw�K���8�'�kN���z9�|>k(y��1��"�-�|5�Ż�ͺ�X~OX�O�G���(�+WJO} ���Y�O�0_�%ʣ��F�XL��'�*�\b��^"�7������|ғv_����1T$��J���Z�-[2���-��7�/7W�ܿ��Tt�ݦbd�
��i؄�B�Ȓ�%����Xm����f��J�hxz���Nt	]=���@���>�X�1`NY/�`vvs;	<�w�S9Վ�N�)G/���檀� ""(w����G�N���۷�R���N�Mz���f��[��uh2��	�!<�����<� �g	��>��5V�=�!�B����Z�6�/����xiM���-%AX/�BL�_�4a�R�����	.�M�.�eZ.g�k��&�kc#A/D��e���ҟ��`���S�H?�y/��5�r���-�n�b\S0Y�E�6pz�9&���g���3��T�2�a�(���)e�W������~�h�dB�Q&���d~cH2�7�QD{��w���-�g��O�w����3+>OJ��,�&W����Z/0	O>z0������������.�a��l�����M���7>�"' ����{e-~���2Ҭ���s��oa�+Q�մI|�xܕ�ꛋ�g� l�^� �i�A)��Ή�D�\����CHw�T�4`�k�P��]r ������5,`Zw/��(�m��8�Z�q�kI�k���9-��i��wor�*%U����v`�4.���$6��i�4����%��5��V"t�f�{
Hl �tɅ;f���.!�~�n�H�a�����M6�3������,�.RB��Y�u���� _��;��6���9��*���Qc԰����~���(=����Q �� g��)���܂�hi�gT��SN03� � ~ey/�
�^�]o���~/�52y�-�{�j���)�?��~3l�3�G����*��Y'՘DrN�k6Ҹ�Yk�2n���b:&K�dK_�=�*
�ǲ������͍ǀSs`3 fk�p�@�QZ���I��E�l��vh1w��T���j��DS2i9>�E����ɇ�-�h��]�a��⡺�j9�g4\�M�<\՞t(xR������v��^� �a��6�h5��ܫNHr�*���b�}:C����͠�~���]B8-��Lk���!t��{�C�N|^ДoU`�����|����	 h�����b�[=�w2��	�9�ՄT�U"S�B�ɧ��6-��uF��`R%��֧����Gvu� o��C�CP(0��~��rZ�Ӷ�rɋ�4�i�h��-�9�k6�		��P�il����a�Řb�0SI�2n<)�ǹ��>�EX�<���B8�h��M@\�b{�(����^�וhGI�ٚb�-Ȏ��4r�ڋ� ������Q�ׁ��]���J�=���8����ըd��?D?��� ����^��� �$TC�Q�foGq�W�?��M��GC�t�� &jBU�f�:��o�/�];��*�D1�g�n�֤h�X���k!G���)I��>��2$^�\8�8d��3\s��2���=�j��w"��,m/���~4��+�� ����N��i3��*>qF�S��S'#��sfC����a(�#$���l�ӯ���a+I���;�M�p�a5�Wz��"*G�����j�^2�%0ɪ��TA���/��u�H���S�4d|�d�{���4�a@��:	D�^��@ඹ��;p��Q[ri%Ƿe��JL	d��e���uz{_���Fr�/�O�u/'���){���8�1AQD���f?!��o�%��p�L�ˋ��s�jv���HS�9��ǽ�7
O��޷��k�!�b��^�} ~6�����Z*n9�����o��1�����B�}��QY�CB���C_D���Ŀ2h�#��\�>4s%%��'��ȻW��3�	�lؗ�O��ڳ
y��e�3IJ+N��m�u
�a������q8�X�E~� ���[�|C��R:-Z e�%�
W�L�����ev���)7�?Y�k��󄲇>Z�UcJ��T�D��E~�֎TGo�z�"�K��&�B�7y��5�)��.J��["Ͽ'/J���`�!T�n�E������2��{���G�y;�G.��k�1?�A룠U	yK�s' ����k��ƿ���;9L�3 y�OdAb��=�t����
�M���Z��>�2���D�?wku\��5�P��<��$�O�].�+pJ�S�?9�G��'��w�Pp4�Z�È�.Id�RG��T|�ܟ�����V��sn7	kҭ�H�I�(����ky���4/т-�as���+C���$��:��]�k��gAJ���C1�>1�.�%��MTh^v�F;��S� ����OKW.��ͣٸ$�^�Dm�V�$۷��J�=I���oG��KwE���" 5T�2��+/j*
Դ3C���T)F�+y�F;'UQ��r�������s��8�����avI�0&��+p�Y0��c���|��q_���<��#����/[<��X�!��"��ƭ��x$=�x����)��G� )Z�K;]W�]%��)��TL�l<y�>w��X���_U�i���nm|wt{Q
��
�\���HQ���/W��D��M�V9;��N��I�T��Ez�{�
���<d��"�B������r�	�����|R���lg�%b�f�cfM�&�	ܗ������ �p?�|2S��]�)��]QbU�Qx��9L�Q�:Ԯv}���MPqnѮ�X��gE��z���#K��O�7�[f!�IVn�/�l+�F���[A�q��ܕ���WPD�PX�����M���I�A����ab	�n9�2.­G��҉+��B/�����Q��R���¼���4)�M��]{�OࡶE�$��?���A�Z����N�\�>�4��ѝ��D����ÖV�%�%�u�LH�K�)������dA���g��a�tuN�� /���3��Dk�D�=�.^�2��� �P���`*�tQÖZ�d����y��;iѳ�g1�0�
^HY-�!���'�L_�0����\��xXF��}���@o]��F��eyNH��*�����m�OK�hE��\<���ӵ���o�LVX�,�κ��':�E����9����!o���G�)�zA��j�u%�����6>_���\G �ќ�6���Ӷ�;�Et��8B�n��c���꽶�]�������]�I���}s�:{�b���Ҽd��U,djT�%v	�����
}[ ����ׂp}���3:f�wu�y[�rrl�����\������W5�dA�0R�%�/�����Sh��1��)��f�)�['��O��r�;��S�RR�<�DE�nȩ�����|(B�j�Y��?<���]�f���s�$Q�h�k\4���dV���_{�
^$��L�S)y��i�|����Ŵ��t�M���Z;A ���^�你�%�ʫG�r?0��g0Q���+��50l3�&�:�L���h83T\x�ttB}�^�������)Q'O7�<��^,��L�UH�=�)Qb0N�6{.�b�����-�x�L<�e$u�b 
鋅��Dx�Ӷ��Q7K̥���j�|��
��$o�iu!U�YW�����[��@��(�0Ձ�6�D<z�鋺&;�O�	G�}Ö���6n����2�;r/��W���Ry���WN���������`l��"����&�H�)��lC4��=e�Zv�?f���{TڶE�Y��dG�;a��h����MK#RuU�����j�(5��4����ta�VLy�4)��=�{j��I|ưA֙�.�jg�﯋ݎ)�� ҂+\B��K�s]����4�Z�?�N��xy8h3���#�0�2�z��Kd���SQ���` 6 �b�&�ۢ[Z��_NNL�)]�s;��QF6,4a5���b+��}㎷�U�Z�ue�{9�w���������@x�lm �T�����@���G'�&Yy�뒚nH��+��^CuNyZִ���#xYlG�&������m ���(�L���j%��:ܣ4(���|�5�y?��k�U-ꦝ�3�|��I/(�g{��߻�X��n�D����J$~@ŷ�PO1�~�s:p�`�;J	!s�ד�Bi�ʘ��93���d�t����h����|���&`>���D�%C4/5Ow�
�|���.����4�UQb����}K��k��L݀G���W���R���p!
:�	(��8w��$�?	�v�2�\�Ji8Kx�M!�{d�Wde�E�@Z�'�5 ��;^��Șh&
���(o,*/j�p�A�]�\�ԋ}1�{U�M��"�0�w�7XM�F�jF,-�Y��l��mJ&��R�n��!p�����F�bh�$��x�/����%O��W4F����� 2:<v$�G�/d�"F����@S-�(_��]d�˸ޤ����y��-<��:�~�!k28��t�PP<l��c!�e�x��-��RFg��/�o�T��<��
��N�nvT��!+L��E~~p>N=6�EU=�TXx��F!�;R�X��O�5�#=��	Y��\�m����m_\$X���� 9ڤ����g�?[(V�y|�,��_�k����T;�4��9��	���Ϝ��;���h�^���pH��9mʑ�2���iV�{ F��0ݺ�ɸ��ݖ��i)� �LJH��N�_���ͧb[��<��a���܅4�:�^��� 3bBx��W��/R3�w;��ծC�!Q�h'wY���.7��Jg��\�S�^�o��X�*vI��F�ua��" $��~C2���=��oޢ|��E���|���J��uAB��lYW�m�śq_l���Ql���9x����ě�ʡ��&��˳,������ b�0���^@z���gW�q{6{�$��O\w�i6:-��~�x��;؆��|6.ñش�W��ӎ����-H0��Ҥ�c�~I�Aז���Z�(2g��:K��N���#��RB�{(A$�-�q�t�c��B30;Y ����E�H�(��`1��`~���y�r}s��C�'�<_�!�G��G����y�x��`A������X>�l��j�?	К6KN�в����	
B�U�E��7����pϾ�I+��'�)�=��q�S�+��3Z�����<v�;�o����V�̬�T�[�������� ���zh�!l����EN`���"�A4=aQ%�g�i/������q*U���Ð�r�\~��7�A� �ek��&|q���p��bd�%�/lSt�Z�/�.w���E�0�e$�^J7�~�ߟ�v�$�	�6��)�Hؘ�6B�+ �Y�N���qs)Va�(�HvP�i��;��״��GӐ����Q;��2ю��?B�����#�N��J�6a)*}��<�8j*+�2iA��~F��Q�Z��r��.w�������M�0�!���K#f}=�9Euo��X�����:�D�������SS�`2��\(�S�n����Ni���m�0!�"�HR�V����{������.��RE82��!}̤c^�0a��;NBy�T/�\����S����WR��R`��������6�<� u o��L��.�O��	 o�29Oɞ1�Y����j���t���7���;�&�F�^�ۙ��Hg��>����+jך��[o�g�l�+�lpA����Z�9��� b���1���鐬����T�0�
��5:Ɂ��ۻ�[r��.�	d��+�h���`����3�����O�\~;v�����d�"rdY֍,�j�Vyz�B�)$���Cw86��O3U���:�M�[��F��'�x��V P����~Q�i(�-�G��~�IM���j�Ք	mCP��H����^�9�F��o�����(��鷥u�"|XC)uԘ�Of��0=�xo�t-x.��_}#��0r�/OP��=鎄D'���_Wb��GSb/�i_?�Ӌ�<5�Ԍ%I���C�<޽�,�`@�MU.3���U��.���h4�6�2�|N��V���A�1whA{Yy�XMW�<�>ςsc+r?���!�@c�)�$QTv���~�1��y7��]�3y聹8����H��^�7��gT��Je���PDr�]���cxb4�#�ʕ�aq�W�@����(2�_�{��$�隣p�ߤ�vIrjuN���T�+�aJ�m���d�AyS�`Ƶ��`^�c�F���T�펶eP�5zx�N��GtE�a�L���2��%�82��jFQ��n0�>�^o k��1���JI�v��Y����@'�7�3����tB�g�bК�ۊ`V�J���2�\@ �b)Mfv0џ�l�8�swE��бI��f�G�/����.����G�4��{dX3�6��=����˔f��K7���͇��W�q&��'Y2��>��*>]�Ldp�o����z���c*3���?^��EMP���5�%�=I��k� af�k�DLH�����rӶ�SR����*U�����A�1��A� ��u� g�fJd�
N+v�-�ș%k�q�MΚH�Ӊ?wp�7C@�� y�9�I�"��c4�I��f��(ZJc�T�"(D��ת��%4��p�aK�]=�nZ��o�Gr9&�7[.�����-�E�-����$;�\�5_;z9�%
�?�c{,�)��0P��3�j�����;�/p���!�=��߱��-_��K�:�A,�K�{��t��H��`�X�u�O*?�|K�@��g$<�b��3I�c<ǌ/��]��y������#�KLФ�J�h-���k���,Z�(h���~Y��|��y������se�P���Ů2�m+7.@H��1t&�Q��|p����eK�3�H����#�M�g��6�I�򌬨��3Cx�C��=�3n�8d9eV���OM���i?����Ǔ��% [�!)2���m��eq�8x��b�;mAב���8��d&��UٺW�yqUL^��.|Հ�u[p��x8�T~�U��V�ֈ@|�}�h~���I�ݢ/�2(��}I�C}ܒ�H[1�D�.7O*��{�?p�Z�:&�;���;����8K��^�vH���]�Z{�_���� �������0�+"�Ɨ��}�����[nK���+�s��T�4�z��&j��(a�ܓ߮��FB��G�rס��nt6�@�w٘���C+*;A}�ތ��~���i��B��(`����hꛠ1tG�y�I��L�H"`�� ��ϓ��ￔh�t5CE������;xLT�p�9?�Xb�1��j_��8�)��/~��p2�/�G�=���*6dcm{89����1�FӴq<ۜ-oBd&���f�}�/��T�9�&W6��r	�����Qw�i��q��f}RRKJ�@j
��C���:ц
Kr�E<g�b�0Ʒa��
Az�q��ҭ����C�����fP�So��?��Ѿ:[<�c�7��4�6U��O�����{2����䃠P	C+y�ɬ��� $��
��㙟	O��p��G�݂��U�% �~���]ʋ����=��ϑ��eI���qZ�&CQ�9��i�D���f?q�XM���;h�U�N}�J�l��?�U���|׉^mFJ�ڙW�����S�{�����>��	�����j߉��Jgu�P�J�t/b*8���6]�PO��$��9uP�������P�HR�i�������}t7�Ǽ���d
Ƚ��DKϲ��6P��n�/�F�S�]�4��?c1r�'���S�q}]�<"62�����m�^��uP��9cxz\����B�I`�!�c�)l���T�f��GU�d��T=݃_���x7<���H2g~�'�ެ�i*��[Y 0�Y�Bᛍ��,�d4�ώ�]&�7����;�l|�O��5�4d� �HBk�[_�%�Wi }x�SY����M�1���w��e�����m��Q�N��r(�u0S��P��#��vyu��o�Ŋ�=>��0g�|wde��D����v��QlQ�Ǯ�c��Qv�D�b)d�멛@���JM-Q���eÞk�!�10B&i�V��$V�ӫ�7�"Ta��O6Ɠ'c9���`d��=U��T����Z5����,-�Y+& �^ ;<����%n��/SP�� ��YY���59�Q#I�����w�q�ݤ�}$@m��p{h�f��	\�Q�aY!H����������\�q��:�	�J8X :�lY޸��Ɠ�~VgP!�:}�w=h?�u�
x��,�lJ;~��uZ�����D�,,z�@��,����Jn��\`A�D���^�H'ehy�v�ik�X�+,�Q�R�P� ��I��n+
��\E�d�M�
���P�)I�1�.���:&�#A���{y!��/��S��Z쟺:g�����FK�I�����^����A�Y��vd�3�:��X�2��+b�r)��O35+��ì�t*�gM��s_v���c��q��.�"����n��12�����
�b�prT�����'JcOh��e� �9���}8<-�	�'B��>���`/ߺ!X��b���pʯ|�wc���-+�*:G��	{�����+��<�#$�z�2�Y��~���G�lOG�f��3���cr�����a��):�1b-G��Pb���璻npH~�2>�K�u�t��e�R�>�B4����~���I�&k����QI�*����,P5��
 ͫ���3�cD�l�|�Zw2A���B���m�.2tGR.�uv�$����6�_#���A]~�r�\�� ��Q��F+�^��#ܾ!2�o��)��3������v�˅ɋ[�+\�'`D�z�|3{m@��@W$l2�T3����[��Lu�:��[4`o�L��%ow�tm�qȔ]�W�y���(M&���v� )p����'���Wߩ�*���Q�Rg��C���'ix���;\ԲMΒ�cD��"s7�o� $7�I��@��0N�i��D�Yܗ��3w��Ny�����P%��!z����h��Ծ�>�"G�M��'U�Jh��������WrF�@?���z8��!�٠z�ܹ� 3������w�T���1�P�x�U�@���#ѿ�Q`gUF��M[�O���+G��]��K
����l`�xGʷ�N�����T�������ڶ���I&�t'��*�W^�/�#����� ����¨�VmS=a@;T^�[�8ŝ��e~ʑ�����0��������d75�r�\d&���b�(2!���u�C˫琷s��bjK=����!�
��Ф#���RS�150��{�CUGx�g��r$$��0$��c9<[׳5,
�#8���?=���Q� -���@��^ʄ\�FA�ԡ�t^�b&Wt����V�W}eo��_���֠xS!p��P�H]~�'&n��[_\)i��uo�Ӎ��
�6�����qdm�=8=�'A�Uёl���!a�d��9��'T�:�w�]%Qg��9���
#K$M��ߥ*>���Ւ*WQc��<T����~ć)p����Hm^�!�0U�<�d2����h��V�tI�	�QH��kB�  /~=U�W��3��Z(U�4�ijW3�ç�cTfB����7"��2xH6 KGV�Cٳ�؞���`1:�`�7���.�i���B�:��'{EQW\���v�q��ݤWM�Z�Hq���Cώff��r3��߇,�jҖG�t��ˈ�8p���w�r�	�Td�ks(Q�I��Q̫,7w�ny������s*l��n��|Y�`��5�w�͐&O�����S4L��mC����6=8�4�d���&�[ۀ��[�+26e2��5#ѵ���M�To����^8RU7�L	��*is�٘�C�(E�M�ç�NX�v�G��D F	���hJ��0�^���&\�5L/����6R3G� 獥�C���-���4jԗ��g�c½��
������������`�-H��zaq�	�ԧ7�A>W��^� Ic�b3^?�Hj5�c��R� �e��k��
�>���x'G7U��o��0�J���n)i�1ہ���Ӿ�.��t���k��H��v�a�
VL�P8z�~��7�.6�~�ʥ�XIR�}h��K�S��E�l	s�Y�Z��]|�6�l��S4�ʎ���Q�Rɞ]Q�v�2\�\Ѵ��b��`��,b��r��������ϋ�a)�P/�?
όݨ�#�k]?t�5
jqת�h<��U�$�֙ �2��%ϋU!�P�s_�;���d߄�����d�?����xEv��Pt6`6��O�,W�e��N[�b҄b5��]*�*�N���T������@0L^��7IUZ�k}o�0/��ş�|쾣ICd:�a��:��4s³z&z���#�����&L��u^&�.J�bLSoZ@��H�����`�K2B勶��b���5��5�X�D�)��C�6|]^�$��.�٦���\��\�p�}_�,���2�0���dO��K��⤜yv�il�^��2V`Z�kԮV�j��(�{/�\�_;��J�ۖ���Y��\"���3gdq{�5� d�ʺr�!�
��0�z�9��sx��;d�_�c7�%&���84�%�O*Xx0�t'M����p��Oۦ��φ��FhetOz��JP��V��I�ga�ܲs��Fv��LH���E%�l�W>À�8�El������PωA�:�K���4�6]"r�
gx��f�ʄ���f3q�����	�h�j�U���O\ �7����E�2~�G<2j�L�-ެ�aue�\�άAgH�(~JQ0�e��Y�d
�/P�B�� ߂ ���*N��W�̷0�ز5���o��u��o�Al��n�:pԳS#���I=�;��d��l�:� k�j�������#΄�����BZ5��0fqf���%ֺ�A�n�;GU��u^S��`�x�8sQ8����_��;���'(g��a��mIOe׷b�����{�c��s/�DN�a�n�z���Ԉ�H�5����i���4�Vħ_��tM�kWZ��7Y=J�7<w+މsK��EroWHr�f_��wb�<Yo�p�:<�M� ��&�R{��Ԧʊ��0"�.X�+1���O,D�%ǿ�Z{����f\����;j&�r��@�` M���kw�D
��_��%v\3����D� �T�B�����OG��N��*B\g�������A��m�p�{o���}F����5�:��%�1O}1���Dw�D�n7��<< �X�b˰Rㅞ�g�ZH����ia5f��ߢ~h5��sL��{#���US%���-�t;uZ@ZU �����%��ʜ�[�T;�	�Ԉ�Y���{��-2U2`���iH�C�n�i ���8�m���)0��ܗ\�g�l'���qP��[�-w����D�r,ǎ�,�{K��5z�u	�~��D�>���D"h�*��jV�.�t�A����~��iO&e0���v�ad����o��	�/p�
�����J-�g��U�M�=)v@�+|�,��k���y	z�+� �o34�O��f���Q<���M�"�&����uC,��#ы����%��kTp��	a��m�|�iG��`I���7o~a��ՅlK�i� {���d���S9�3p.��%X#=��2R�ke2��b�Ă��8a\Xlz[A�h�\�f���0�x�u��Q��cq,�A�g������$;,�ys�Q��O�9V�"�͇�+��LtAD�w �J��bf�* ]iQe�j]�j�0��ſ_��5���o �E��*��������U��mx�b�O�'v5S9�l��l��2ʧ0�d2'���:Ѭk��?R�2�Z��B�F�|�朚42���Fk�d֤�J��@1�M��ܪ��%v6$������R��O�c�+-}��:� ����f�S*���VV�R��,&��4���!�L=���()X�P��N��ӆ��r��k4���O��#��U-���i�.��s�֯[�&Ǫ̉��u��]���W�F�B�z�hA��qvp����J?�{�O�/~e���r}�~K�d���i���ďf���)ǀ�ֽ^��� M������Z[4p��1o߹S~ ��2�D�f�>�r�d`�Py㔉SAD7���=��fuJ�����%I��Z��O�\���OY=��3�dw֞\�p���.��T�kޗ�L���ɶ��G���5��"n������!$�����M�e�a��O?���3��"C��U��%�������4u&��X
t�~��_q���Z�:  �4|kPr�J��Y(*`uEAiy@
�6�3��˼�d� ��lZ�C��<ÉW�����@��d��P.C���7�7�3"�R��~ժ`��L��"�qۈ��
v=E�N[�@m����T�7rۯy!�L)�e*�ż;q�r|� l���_�9�9h�`� I���.��J��L ��3�w��z��&NHG�+��?o?^�g�>���;���C_��lm�ƆZT������V�P H��V��W@s�`r�!'�F3a!PڮL��-��In�L&��=w'���nUκ	��^���!'����9�[���d�ă`�?��[�1�7���-u�vK�?���q�J��I���ݣ5T�0[m�K��G�{U�����d�R<�b`M�����Y��u��_��P�I�v�g�j[��t^U�6V��dB�K���Y�s��c����Rq���Ҫ�׋磨�a��Kw� |��4+"�n+_l
���~k5a��F<�!�
Y�>B��������:(�p�m�O
e��9ȭ�r�����|��B$=Mg
g7����-VZ�x� �|�n4���TI���(�_CWm��8=�2���D��o���j�}�P��wf�G
�(�U����^��ޗ�ʶp��I�JA��U[G�q�=p��v�����m���)ۓ�x�`e��7�]H<^�uA�bs��5m�n�_����H�ɲQt{��A9��v��~�2�ta;w�üF�������;y���,�'�Sp�[Vk'a]�q�Tʷ[,��n�Nc�bk��`t,��j{u�M��B�����</#7+ 
��D� ��xQ� %Yo�
8	|��rdR�/��bD��L<U�@���H���&T�Iv�����f������Ҟ�跟�d]|t��	��[�>��.�&&Ra����� _W�C�b���?7>����[�iFe�C!���a��]=���T��R#,}x&�����.jb4�-Yl�����Q�P��WZ��\z���VM{5vTK+���o��^�݌/\_��~y�	��l��zm�8+{{��H�4��.�幘����\�R�������PCnD�2 !�m����c���`K�n�6�"���]C �0k��j_���^D��) w�0��ʋ�՜(2���^|����؜2K�s-*�����-���unx��'�ˣ8Dx;�V,$��h���Ei��r�M;�WSʻ�b�#W�DɄ>��h����z`3A1`I�l�����������/5[�0�ķ��-Eг���e��ϛ��������"��2���������b�z�}��|�ɳk���A�K�m͹�J�T
�	+M�H�̃�Ƴ�&�!��Xm�^����f�@���(��-��M����Hi�g��u��/� �C�jxn|澲ا��<�{:	_gX
s���)�����
Q�	-�O{p���<�Na�1�:%`��I�i���'�K��ʩM�voa��/v��p�|!{�CA<�rR�訚��mY�6�Z�!�����We�����=՘7�U��ɵ�SEB!���|�j3�vu�c��������8#���R�V�����|o��`�N���E�%����:���P:�'��@�, '\�~΀k���i\�!��B��X:��D���s�w��N !�nM����1�Wq\�u�w�M���/4�ؗH*v�������*HC��̊0��x���B���gBF���^&���˒��PY	�Շ���,�K���'}B������ [�^�����dy����߆1��K��`@�o��;��Z0�)sR-�j'+�w��#��>�L��)]���]�@$�_�-��g�'k(�P��X����T��
��x�uAr�$��d���w;���D<�MxL��\u2f)Ӝhi��7M��^�J�R-�-��y����!̈H����t�=��;��:�Ā��ƮU)7X.{=I>s����+WC��Kd�m����h驴�Rx������#~`�b��#q���x��%�B�7��Y�%&O
��*ɼ�D>ㅩ�3�M
�Rٓ���x0��0,R��w��+|�g	ѣ=9��Y�6��/0-LF]�	و���k&9��al�m���d6~�>R�0~l=go]B�Rf��*��V�x�N��+�y�)��p1 �a��'���4������7�[���o.�"<�l�%/�Aǆw���`�Q����M�����a�N�q��F��0�Q���
�{P(3w)k$��׾kI�G�(�M�!��đi� #Gg?�S~�OGf��B�r� !�&/0��qS��Ņ
D�_�Lk��~''�;	���@���F��uH��W{�VǺ�Y�5ӡT� Wmސ��2K����
[�#�����E���@�����WSd����s�9���UWzg[Փ��iRZ��&�k�P��	� �F޴��{j�Z�@���7&Z	�����q�7#��nF���
1@�g�G����n��V�	ݮ�
����=Vck���Fۉ�� CQr=���c�U��&��:�y�l��Rz>B��6�4m�mSc������"���ȂF��3%z�lN�>$] ���$���`*O5e8��[mj�#��_-�O-�}�j
p.zȮt:�E񘚦c�?��ǐe��ġ��\@��͗i�f���kKfQ���GO2[�^'����e����:jObbיYU%t�iq39,�1aILB�b*Ӵ��8�����"z3ݶQ~�}�	�1 Z�� �B1��F(�_1
o��HIw0�<"�3��9��O���v�l��q>{8f�6HFl�]�i�R�| a�z�#`\8��23p����R�i��vC׋@�����&g��_�?��M�-̺�z�sB3���#�ҧ�"10o6�{ʖ�-���w��E��9�Rߖ��`:�#�հe[E�?�SP��|!$t/�*vL����T��fW���vmD���iuqY+d���͠��Ę>×��$jڬ���q`��廪5K����Y����Q��ъT�qWl}:xw�b�r�f��t	����d-AV:��@�*� '�5}�)���0��FA��5�"��`f���V�F��a<p�\�a ��x��r�� ����3\˳�����r%Q�kt�QX�0�q�R��>�d�]/�6�Ò!�Ʌ�#.i���u_������Ŧ;�Q�?1'�1�zrJ��cz����vvd)P*J�ՇB�����0pȟ�p����N'�(Z$"�����d���sFx�e<��cbr^*k��wFOD\�sㅩ]\Rnӽ s- ��,�wF��+��'���Ͷ�hq$���H���z��M��1d�f�#g Q	������Y�"�$�xK{U���û�J�x5,�s�U���QAd�n�X�T'�V&�	�'���Ѓ� �?�����H�>���mJ"���J�	�p�D9-�&��H�м�lW(�lh� ��~��9j�w�5��m���P;�z����hk���#B�o�u�Qh�xe����x�RRe��]��y�N�0��X�8)@��.��B��/��K�!��s%jO�0z�F�@�-����թj�֨�`����P�R���K�������,�jUr� ���+��:� {��y� 9b��Iv�1�F
��sq��̸�_q:��
n���{�j,d{�j��}�h�����c��ȼK��ڜ����^b6sh��dN��6L�#�ag��N �ɺ�/%67"~�ڦ��mM�6�'�&��������A:7�q���F����j��v�=ɷBzH`�*��z�0�)�]Դ��.�nd�fJo8`3�6c�T����}�6�UX�r�iNv�߈�֔=/Cf	U�sY˚�t`���� ����Qi���˛3�5�Ý��c-��L�6d��B]��(����A�c)R���VC���;w�P��QSc��``�u�'Nժ
G�v??LU�{x\�N&Z�شO�r]�<Ew��#���y��zq<Nt������ɴ�ψE���՚�K,̬c�}JVjhjfu�(:A$��p�!�7�C���&���$3{��G���)l�x%�(.��t�}��o3�O\���˜s�f&B܅@��}ث9��a�^C�:`oYn�مy�`��f<Jz�X�����{ꃺ��`afw3��&k�gL�~ߞ�(��yG��&��SPY���r�r�vq�	tv�[�K��d[mL؛Ǆ4�NK��a�g���hFu��� �DY��:)͹�2KG��g�
��D���K�-���L�]�=��H����>s���d߀���������'|�a�I8"����g���}$�[u<���ۖ0&���}��y�p�]�L��ŧצ�Ub������s����)��|B����\��y����g��� 6`�HD�XZ�>Ŭ*z��0c��p��R�M��X��?�Dc"AI�V�F^C�H��\�k�@��8u�U9eq�q�ڹ���%��S�܎T�i�[#�yћ$�2������]/An�qp����I��`Mq�9�� nT7��}�}?���Тn��'i'�h3K���|��*\��	����8�c�¹�ѡ[
a����������<%̇N�:^�")�c�R�)I:�n� O�oS$џ�Y�j܅�m[��Ii�G�C�gJ<�Z��u�ޫ�����jxd$06�
:D`�>)/e��BҖ�~�_k�q�v��>�4�ABO��q�<W��a�#��o���_k��ڪ,��h�bWm���1�[v��8�7(���}�tx���퓰K�eTLX��/n�6�]���EZ.�o6�Wq Ͻp�"���+臒k�o�;�=nRW�^����e�o���~���# �0_��/G�Iea���=˞��*$-����/-IZn��i�R����v������=ϱ�y�����xx.�Q���8���]��`$�ۆp�L(�+0'�d�L�pؕ��6��D�c��To�Q�e��vw<yY�zEX��J��l�2�?��t�<�N���������ߦ'��$�� nxm�{ҥi�|p�,����-Rm��_�������7���a��|���i+��Ɛ��ۋ� �=H�(�췲G\�)�L`��*n[F�.���`/����b�P��tP�V�l�=Nșh)5TEO�=6��!lg�G]�<��MQz��p<_c��Nܚq�7��ңkj�B�ԭ�d�+��	� ��<��~jh���o@��],��D���T=����~(f���㗲��v�ݱ�RS���-��e~%N�/���e��/Z�,��\���#��j���ǵ�z�(�5]ԓ�.x��ൂ�4��+�g|�l����[��F�.
�J���b�6�ؕ�C.�*I��+�๖tS�Y9��w` ��˄j��g��I�ˇT
���mދ�ڍ+����S�x��J�	(����N����~��_���>NF��n��ļk8��
�Q�3D!��]i�6H��d���*{��pr=l�~�%)�S����3������`D��	���uU�����@�G�"*�-�aa���m���sɶ[~β���4�=YF�>֌�9h���-�z�GvZ�1r[m:��8����$��;�3��2���L&��dҦ�af���A�[����)�&�\��锻�gƙV��oW�FDֵ�Dj�u?�l��y`s�9��a�43�f9c��(��j�ۭDU���WC���s����?!���*�����:�ޥ ����; Os�1ACg�frtZ�l��:������p�������Tc�7m��O�	l��������r�5�`�J����P��C�^�9���$� ʞ��T,\�����Θc�N���c{v��j����C	$.A.[��(�3��@)��p�$$�q�g
�ZV(x���U�z���o?2i=�M�b�HӘ2�D��E�}8���[Q_�� b�TId�dv8�\{���am�c��hz ��p@���R�@���]3���`���L@�n���ق�<��#���Ͽ�8�øwn'�m�L��-b�vzF�h:�(��rY:�W��3����-�����et���2	����^Z�U�g~TKBfw0ʓ/�W]2�Q�	� �,�S�}̭@��d1 ,��;9oo���>�����G{h��f�5TU�ԥ���Me���e�Ly��!�
87��,0:淳���X�掫d=��X͠�v���C��J��Ŧbg�M�#A(m�]�R :.hl�a�l��#�y�	�}�0�I��f8ض�����e�f2�l�e2�c�<�K�&�/\hՏl{�g�7��i��`��{���ԥ�5MbΫ��B{L��#�|��(�@\P)�1!<��b}B���2Q��ˮ��G_�:��P�.��%
�%F�$UV�wO3��v!�Yp���&�|ԬmH�=պ��eؕ�Uˈ����[;0J�'�c�O�$��W%N(o�2wxW�dsB6/.��
�P [d�C��J��X�c9K�*V�k���e���׹(��B"�j�Q_�{�>J/��P�'����E�9����e�R�h�����R�-�x�&�� ��;�d�r.��~Pl��ɂ3Ww��=�Wo�zd����B;Ba3�҅ 關WbjYD
��,�s��-�`3G����$��г�?sP��Č�Y?�sCK
���`ᛮ^A���j�n�[����x�,��<�~-n�Ut(��u���!���@�t��WI&h�uh�;|�ך@�=�;�6�&E����,5U�O�'�� ��Mx����ԅ��ˈ�C��r��< �/<�PaY� ��x�F$������
9��؎�ru��:�
�۹D�m��Ơd~�m&�<�^$�GƢb�� ����M�����1�/_��MGgk�|ޭ���Aj�g��c�H`�N��:V����ܩ�(,�6f5�L����j=��ѝ"j�!�M�奠}��[d)�������є�Y�Dr,~ߦ�Z�XZ#b�E�Ë�a�Q�Q8���ZV���F����]�2����0ضe�����T�����.��O;�@�� �jw�;��|/���@G��c�h������vJeԞ��-���rrL-2�'�n��E9�1�uQ�D׻��#o��m�X=�5Y��r=��)���-�:j����N�زbL��Ѭ�n��Ƃ*�X5̌�O �ءd=�O;�	X8=@��6�\-l���Sh![�������z�Sr��6l����?G�e�g��{%_��.����Ѓ���)9#R�&��bH�Ӟ  AU6�)����o`�������LCjz/s��ON|�H-��D�I����](� m�d:��BP�10r���s=�烈@�j��\<���ɬ[��z�nEN��h�<�
\R�����c�܄���m�/�����r�uJ��7��TX�b�-��$>�+'���9�U��V.7�(9��p�~��lo'�=B���GK���dm���f���:�:z*�����ޔlO|����2���� ���Fd��������iI��^����y��T���;Ҫ� Ɏ9�����Y��	\��Ğe�B#��BT/�0G���Q������}w�ў#�ZMsvα�BfT_�1磉�j�j��̹�t\c�\8A=f��]&7ɜT�Q^��A�S�|�7��v��Z<��T�T�V&��x�X�@%�0����ԕ%�W>�A9�k.s��)K�%�<v���D~匍5�P�Ҡ�`^35YR����},�k4�=���q�r��j�}-���l�}Q�w8�cD�rJ�,'�d�ټ~���֒P:��-�Zw�W�&Ⱦ�z��]�@�~�F臏6cPw$���d�?·�@d '�q�r��L1c�k���׎�����aX���!}.-W�PȊ[$��������<X�iH�sI�p�b�:��VX���b�i���L��d6O��keN���,��?�}�Y�kt�HB$��UU�s#��>⅛	���;��I��]XO)��l͸0������A�Ͱ(#�c`��aX|�_��{!������IpE�R�K��;u���f�Ya2���wC7忒o�vy��Uw~�)ƈEc�d"�����2�w~�;��$�Ĉ��ԋ����:#��nl�Xd�@���*ghP�<~1غ��?��6e�]w�����W7�#����qk xi|9�ZG�R}��X�£'�g���ʲ,�$����X��y	˓.��J�xdV���u����?�(��Q�!��|����^���
J�	���v�?a��q�-��H׾"�v�a��M�x�{\W�Ŭ=G>;�}��I;���!��nWn{���و+�#3�P����3��y����'ědz�� Ka�&g��<������!�G]|0���D����t�ڒQ�߰B��T��+sbr�D���SݛT�JP����C��	��T ��!n,ϊ	0V�C��P�ǵ���劣!2��͐M�ؒ�d[s������m�K�t��_��3Y���B��pan��C=��ra�O���ڊ�Sͫ�H���Ѣh���`���ﺮ��Y��Ld��J�����:�+cD!��Xdssx�=��]�y�"�X�o�q�*J7A�WIw��Y˾�nT����8&o����l�,9c���trKREQ�K�){R��D���>L<��M40��_�[��#sR�w`݅���Hw����h���x� �~)����4Ԣe}�~#]����-#�g1ab��K�|	8;��vq*�04 ������t���c��m>}��aAR��B�t��e��� �1���͊e���ڌdè�4y�+%���9�=���j���A7�l���w`����U󧼤@�ጣ��ߓ� F�'��WZx@��0-,k�����w@���*��~	T~7�h4^�O��}k�O~��S[_�J{sa���q�R>'�u�n����=��u���'@%*�p���·�H���9a ���s.\sM3}��L������s�f�r�?���խ66莡�F�*�6c��UV���r�҂�P�ߊns�}5�?��Z�+�x��$�p�Uƹ!��հƇ�ɨ�Ա��/�jt&h?gY5jR:�a6�yz@� ��𽿑��A��i���P�A�:�&����s�N�ѧ���5�2��[�������2�J�1g�i.���[�%�a;��]��=a]���b�W�[�	(v"wv���f*UJ�9��»��w2���Cy?���Xw�Gq�-��6��S����J����l�b���b�XjTqhۋ
@�^�E�M��~s�:��`����sIX7 @�@Ӿ��хP�J�4�.�h?�"�_UO��($��ʜ;��q�F
���1
�j�fn��������x>fN�C��:`�����_�1N�Vo������v�o8�[^��%L��8Ȝ�1{�N��ڰ�S5{�R{���i���}-�s�#w�L ����e-��� ���ӎ�5�F��s�� ����40�@�넭ijRwQ�?zf��uPV�NA�*_l�B��m97��C}-�l�N��"˽�k��uݐ۸���<�c;�ۿ��Q���N������5�G�`�'CQ��@�0F-}����sl�������'7z�gZ������E��/#E�������U���c�-0�f�G-��t�祆�Bm�Bj1V�Nh�RAu�_�3��Գ��� M^��v��ض1�p�G	�OlS���-\+�}���vh/���ĹR�^�%�[A��Y�� ��ZUK��/�"���ZfZ�X�'�B�3�E�ב��[pQr8n1���Tu�4dj��*�2]��Bw�7U�s�tE� ��0�6����^������G�3_&�\ 3uxI���"����!P�X��'	��`,@�^����+]�vT��F��s�@�]]x��=�Ք����Աl������x"�u�3���Q��,���E��T�yoH��ͱ�q���֩�^T��@��Yfe��Ǿ�$���T2����Ke\�6/�Z�:�(}Z�6!�}�J��/�G&c;�8ٌ15TR�쯌�y����%U4����_m��[����X*�D۰�E1w�m�3.��>�٥8���zO=�����ľ�[�.�+�K��_��!T!O��g%�w���^w�v�\D���1���P#K+�,Z�N�B:����l��d��ެ3��Rf`�$��u'����~���>C"�il�K�h;'����D�^�4�կ��б��%?gɕ��ki���� qm�="DKpO���p\US��T7���Kb�%窲^~͈v&O���m����=�<&t����sWm>���Ok�D���n����X���331���?�e���)EvCE^�U�c��J�y�s"S9ְ��Q$U�) H�{޻4���� �9qsm��E���ia�>��W�10��Ao�k �רXS]��)~��$v���/�݌s��;S
��V�od�4Djr���1
������Ad�%?�O���͗�5N-�&����A_�O2;PX<깸�"Fv�VPdJ�b�O5h����Fo6��蛝�|���]��� �N7I2���X��\����q�oi*�3y�s�Wۧ�{'<�Ҙ�3õ����dq�<�w*��MI�E�t1�v�AFZM^�Y�8��b�K��B�嬌�!K#�h�C6��bM�؂Y_]��.>�jL�M�^�F���I��E3�[D>0E*>��������"o��p�XȒ��jc�[g�p�ߛ������9|�Z"c�	&K},��2��-�y@� C��ފ�HpY�	5�K*��	n& M���Wi�Tq�����@<�!:>:�+ǂ�Ӊi0�W�Jz|����d�Yb�=�Il���q>��P1	y��n��c�v�Ň��|���x{�w�p"R~�!�2Y?�$9�qvz�A�r���p�}(f��C����]=<C��
X��>�/z��KalEnj��T�d��=���&_J�.�b��$#��[���Sv���5s '�ҵ�E�	�"b7���?�4Z������ڏ�CI$<�t@�̗_6-�7)Y��(Z~��;A�fo�<�w����~�7�|��/q��Լ�� �:����8z ��$�>�V��iY��=}�k��=���/�U��O�e?W(��Z��ʸ��[���Iz����� ��������URŰ�\N���4���?��v�l���Oz}aԀ��"*)�TCZ�+�����#򎹐`_2|�p"�3N�F�x��O�������d�蝹ajbLA��y�	��Y���*xֱ(��BkZm.��ư��-P��4��Wn%�O��#�mP�2�ۑ�'����A{������|.	_�%20�M
���AvQ�t�����t�2ޟ��X9��-SdC�
A�7�v��!AQ����^I�B$�Ұg��fe9���cL"�Mm�� Y��=��I]�+�2�ݓ�o�y-�<W�$��]�t�d;�T�ɫ�2�kИ�.��d:P��6��s�^Mudmx��fU�٦���(}�s�h������ �yN�U2Ҍ������e�:��Z@h�+�,���c����@V4;I\�&��̰�T�q8=��C��f�{"��VS���'�4ѱ�'�/r��A��䠂�k~<`s����0�*{Vb�	t��ظ�?���R�}�\�Ax,�����ː��7�G��ݰ��G;��U����/
��)�>C��?���$B�*����W�y8�)@`�^�+q>Ν����?;�9����M}�O�6T�ٴ1"r�&􄃻��	QX2�R�UR�V
��i�J��7:@�����܃��i<mL�n�oo`]�ҏ�1��#B�zE}��B�%'�넀��P�����^�B�ʸ�vR�5��y73��k�9x��M�.\��@'�o3�@�8�v�@����|�p>�h��"[��q�0��4<�<qP0�}��pM����c9�o�6al�e$K̑��0[�,>t�1d$%�(�����`��9��}�}n֭ ��Q�gz4��5��^ �����h�]b���Γ�>���<���-[����ʰt�Hp[�0J�lB`�6G鰻��L��. {W����`�"&��3 ���ӣ�ш���O�Z�?�.1�ҕ�Pk�8�c�1�YT@P��'e���R�����8>GiEjP{���x%l�A�����!r�0H�¦ڌq4�Ku�+���m��(`��d�|��ݯ�f1Tj��z�4,[=��
���7^�!-%C�����~
JE����
G�L`����۝�(�S*��G�.��amo��o�	�s#���<�u}���R�$;�$	�z���{&.����"(IZ���6��ǩ=��A�]�%p1�8�o���Ө*���x]M�K�����jܳ��ԫC�\k�d���S�8?���=��攙L�O��)WLs����:�����3,Zp  V�VQ��Ch�L6�R�����|��z��f��jp�3ϢOy�����$X�����$�N+;��ϸ8����È.Ҙ�ފQ9�D�J�/
w(��J�M��2Y�DK�|�+Xl�����3n
�ۣM` =���'� �(%>�<�:Q�a������ci�H9�"��>Q�(�d\K���o��v P~1[��f��@��csܒ�&f��$��tX��Rq�*I��Sɫx����X��p��؏���ދ�	`	I������,cH�v���/mB���ܯ�hK���:�H)�F��>@� %@JV�j�15��*[�7&��lj�{k����:�oNE��M�a!�_��#l�3a]�#P/�y����}�\�����(�����<hsV@J���{,.��������F�.)K��Nsu�$���|�O:���>�`>�_ �C�������A���N��NZ�fhQ �Ld,�3�~b:Z�A��a"���z���޾�a왨�.��� V�p�%��!��1��|�\4�PEc�wA@�"���%���~��UezHğ�^4�p��w�� ��Aq_e�M�?JQUk\�,ϙ�������^N������l}�B�mἝ�<-�>#�J >���KYs��1�.������q�,!?֭��Q�w���7�rV�L��H���ɘ��F�o��22�z@��`D�� 0O_��Q�ј��y��݅�Zc:���OH�&�Z�BΒέxr�Q�<��4��c���=�f�����oV�}$E#r�qr��u�C0YC�/ַ�Ĵ+�=�j�X#�\�ScT|Mr��I%ZA{��a�	���_Do��>d l.]\�*m�$f��N��Z U���U@ph�+3�j�"g��׈��!�&�R!���@H^Qͩ
j�-^�N5��tL�������һV���e��gU�Sx���@8��q:���螚}���P�	�<���vCn&Z�9���<�6�J��|���`��_�O�q�j$T5x";��g$,�=�*����'���V��Ӯvc�C*?*�j<�v�-/x���u���S{i��V߹ۊ�3&���zj��æ�Ŵ.`�l��/��a1ew�C�D	 ��Q9�w65��̓�8�r��rΨ<%��B���
R4�����<
;T��c, m̆>��|&x�+3���ea�*�EUKk7h5&�	�;���]<�3�dl���EN�t{��:6�Ъ$�
W���+�)dZ��r�N�t ����ň|l��M�s�kUE8�QP䪡T���e���{sXd���	#�X �g�ͪ��ON�`P�C�v���*m�P�
i'I���A�|�  |^�pQ��,��]����$3��@��_�(�A[�p�p��ȭ���M/�������,���ǳX�r�B��B	(g=�:g�m@V���]y���վ�G;E|��v�������B�;7�08,S
D�����$�؈âlWI�9�3��d�Fam({�R �T,;�ݏ���f|W��4��?b��.���aE��l��S'��"����K��& �̲�i��{����*��}�����1b�LLV��kԝ����o�� ��mAȫrL֎Z����)T�Rr�����;�trp�64+5);�����n��*W޲�l��.��2I�"��v�"�������%B�g�@ d��V���J��Su�mz���k�Lh���NHk�_����kimO��D�\Dz��s�M �I	�n�5�OP$[�SzٚPi�:�1�o8t:d�p�q%����V�4��d�u����ؗ"�m�t�s��A3O��ߙb��3�n�gN�/b4sW�V�z�4=�8�+���E*�� ESky��oqсO ��� �gRDh~O�'/��'�Ɣ��'Ӥ��ս���'i�c~g�Z�o�7U��aѯ�C�N��*G��Qjx�1�.���'	�=2��͡b�H�@w�1�<�m���Jǵ-�\������k|�O�4��-��7yz��^�(�A(ڄ<4A�>�K��h�����{�h[Mș �	T��P�-�H1���]rw��ǋ����>8��ą�%s)�h����Ɋ$l�Dr���ԑR%6����Kc�N�ҧð��Oo�9�k�kUz�yY��}@�ཫ�Q�����D��?C [��3����*BJ*Ä�b֞u�픗���#8w<�p,-��}
���t)�lf��J����o�o�d��i�5���nշl��6+�b�8f�
�_���?���/ d�$�� xF���BEY��J1p�w�K%|R)O t���RIma������n��M R���@Ú�;
�^��)z��1! \)��˄Մ����;|Vא��r�1��--v0��4ދ��zt�2�0�s����:-�}�Y��UO���ꍄN��~�ͣ�+�A���{f���C��k<RnY@O�	@^���lh"F�"�TP�:��h��.�+���:y��1bu�N"a�H�f���*�L�i��ꓥy�9�,�:���F՞>��:ebg��n��۳R�� Ւ\a���nGBE�J
d�D���?�{��Y�ZV�F�K�1�7405_����<6[FFߧ�J���T��O�1�\T7@]��7��Ԁ[�����dN�
�b�{��Q������j+'; �i�Ψ7���F�\�>,�|�5?��� &��RW3�.G����2�:�a��}ޙ�[��d1c��!ہ�!��C��O�	�(���Y0>�$��M�x7��,NoH~CNnT:��1���;\�*�KRLp�UY���aJE�?�0z�L��!�Z ;<�V�3�[����n�ˈz �DV��'h��be�3niChR�D��V���י���D8h�"g����SV$q�-�� <B��PƇ8�T7#� !�2B+�)cSR�v��M=(���u���GC6�������P������oP-F[������<av�H0'H�^�o�.>�~�ոx8��ϧ�D��,+�B:B��+����?��*������!�!�v��R���.-ƀ��e��G�/C�1��`J��œN7�N��<��\����D{B��������G���A���Ű�4����b�+�b8f	�1��+w煵���P��5q1Ȏ�v��&ޢ@F��7��ّ����.ŷP\u8�s��� &mf$�-�'��) MY[�4�&��	�k�h����G�$}ԧ7�E���Wڈ ��;�;�ԃ�F#^f����<.��iO@]��������m`�S��ǜ��@��
rj���L3�f�6�w�cz�P�1]>a�q�j�M<Z�/qh��� �,D�
}�n��d� $`{ݬ'h��}�ZrR��������8h�����ӗ�7^�aY��B��C��&Χ�30 ;+����k�A���L�Vd��`��0�Y�R`�!v) ������:T�8*2�N�+�xP�Ļd�aە��aTRY�!�ܼ��9~4F�-���gǧ�R��u�ûv����mg���!ݠ�+U#c(v)i��z���.��� ;�Wۗ]:'�$LG�fbv�e�>#3&53���3g��lU��ߴ�g�d#g$z�u��l4�W�9�&�aY}w�\&1,�&�x�z��~��u��)�6��P�JM�;)���Ñw�Ste�����Adqԗ���B�s�P��h����w��,�S�U^�'�ѵ�2S-�q��S�,����a�D��pG~t�?��^������4���܂��k��dݡ�>�-Ҏᝢ ��lAЃmh;��	��TQ
���ѫJ��b��y�r+�7��g���(�nb����
^t�� ,��W!�v�~E��yq�E�#J�R���0�*�F1]AV��[��ԟDWs�W*X_�ͽd�[�s��c���|.�:9����c�P��_N��1��$0�K%0
��$��>�6=�m�r ���<�sn�(��/���z�Hd�60�:��tB]�>�t}0��V2܎����	�ގP�k��o�� F�7 ���%����.-n�u���_�;+��w���»�ǰ�Y]l�{\Wn8��t�����f7Dt@{uzWN�����'Y�ԯV�*��-�O^}� �{e�a��xg@Z}^&N>@�����2�{�P|y���\�2%��H|Ԑ5����ח�;���h�E���{kJ�����ur$M��
0��ټ����&���u�ב�ވ�}�������8���!
��h�=`)*U����c���=n�攫\`�' ��8�{��G<ˡ�@	 (�hϬm��s��(@��%�2�w7�Wj�.ޤad��Ώ�q��]����/�g4!3$���$�<s���ܝ�Is�\��m��J%�s�cR����D蓀���#�����љ�݀!��4�h���[G���n�}�K iP0/�)���t�,�E��/a�Xq8F���p��y+���������4�
���a9(����aO�'I�Dw˕ڎ�_���]p|�ϭ����x������N��u��x�
��.f@W�A`N������§6�������߷%L�w�@�:�霁E`���5}[ҭ˩�9�J�2��
k}WrbA��Z�Qۡ%����V#�l j�l�k�Gڔ!p��ނ��p7_{W5ʞ��;�{[#|Q�g��f�5�`��B�dD�}��* g l���Y��w�HFܧ���X�Ƽ����X�4<���aT�4�J��AèZ$x����ΡiT\F�
|G�d��%���gz������k�;�:��7~��i�|��LIwȥ�H�'�;J��n62�If�jd�SG��4y�Ș��~�n9fi��G�D�$��b��^�XP7;�ék���ѭ�� �O?vI�T��T���,�`�\�kK��㠪��;U��4��v뗽�	=
!d@wU!�Q�)�20p�<X�玍�\Z�n{ҕʾv\w�%��8��[i��?zHL}�
+��j]xsyG�\���O\��R#6{>/���k��c�N���)
�37���=�l���!�5Wu���R�����9���lĿ9/� �@yJ)��U2-��<��w�AN}$M��ؽ���^�&�0��t�R���(��)����ǺМu���=�[��-o�7�g��8�>�h�e��@�Py�>w}S��CFo��e����÷V��[G!�c�z=b>�#��"g������[���u�����{�ɖҨ�m,�=�}Hѷ�����J 1�aŞ�K�ԏm�L�K�aj8�x�i�{0�mX���F��TGS<k��Z�T��J���'/���Y��ƍ���"`h��k�mJ�RB��������2�g4����=�XlcZ���iR� zk�����ě0DP" ��
o�'�v��or���� $R��C��=M��	���Vͳ�˒b�w7ڼ>H� ��gt�3K�l��oқ�ɤn�oA�B�+����J4M��
#l�]ρw����Pc}��������=y�V�ص�*2�-`/J~]X����\n8��<hb��l��A����0��Je]�{��
>�Z0*S���~YUl.?7�3�1שּׂ��Һy��K���Z�!��q�\�E��8*l� _e����< ���I �w>G�� �QA����Ǘ������m��h�a����{˲���O�+� �{Vm�@&��l6
�z0-����na���h>5`�S2�ڇCx.��Fu�uͣϔO���|y��Iܚ0^4�Ne��\ӨuD�Aœ-��[���6��w�̺o¨������f����}�$-:d�ְ���]���krJ�+Ǩ�%�����~y��V�۵����',s�"��1�͋	������z�)˙!�#�[�~���ƌSN�~�m}���:x�Ԥ�k��]wŽ��D1�Z���W�^�bkn4�:�C�l�
�\Bk���������&�ƥ���gj��sk;dS�Dw�Ϡ�wM��0:��kAuO��\fVq�(A��V��B=S�C�z����{˼��i��r|��E��d�\ng�D��(�NI<G�B�+o`���A��$�n��%��i[��i�܁++�y�t]b��t��3m>���Zv-G��
Uس8���gvB{˚����D1�m����Ca$���*
%�����D��ۿFj�m+�םUX"����	8�<KХR���1����!�6�+���)���Q%�L�$��_vP���|#�4�U�WE+vq�I��X�@W;�k���E�ێ�ϲ0�%-��c@�_i�X��m�����[��6�ks	,�p`$��A	��x��ĺT�lu/[:�4�>��k��9G�i�O{�V�Bl,���&I,V�>
:;����u[�o{��������L�xs���k�6�,U�>�Zu��q,\��L[�ڠ�i���5�n�LC�B-9+�q��z��AN۞T�gY�Hn������<��e�N*�],�?�)���mv����l 0��|l�}S�x1�o��a}��ɨ�ek$��{q�����"_��j���".�ő��5�S�
�vt���k�1xP�>:[
�e	S|�s\�3ǌ.����6��T`��ˆx��H����&
i�2'E1hLk<]8,���c�oLYS<���i��R�Y����m�d���*;��$�Fk�L��p�w������Ҵ@L+H��7c ���;ui��-�6:�ʐғ�̎�~]�věY�(Dn���i@b�)6?�����>$�w�a,�N@"cځ<]^�UB�bF�P
yߞ��"��� ӑ����N�X��\�#����}crx���C�I�M��[V�u.Y��{k/'����]��%^�|�T\�YW��d�����t��P�ZGƲ�e݅������+ ^�d<��d�x��!�D�<����l�#̘8���b�9\kAU\���>������eC�R��s��[�T=��7�ȩ���ʻ�PA��a �X�p*�D"����	4��;�!��hdC�e�#W"g��.��_�Pbu�a���ɓ�JF����y�Z�|\�d3� �ڿ^ƟM�>͔���=S���S./4"6^5ߧ���ɻ�M��������z<+)�Fm�@�6b,W���]��65B���Y�Nn�qH�~/�:dI��S���гNR�b��9Qf*�l�$}�1���0~W��.f�D� ���D_���|9�CE����fkVx����②L�l	Ai��^����J߶�Q��sw
���D[�
R	F�q>:����n�Ѐ�K6������$D�u����K����_�����S���s�:�F7A�r*}����LʍW,�j����n�'gYX��F ~�[ǁ�3��y3_Fa��m
�t��n9��G)��D��K<3u��86L��}3��.xƒ܍�xJؤ�e�����t!�Ӱ+��vg���b�Jd3)l��қ��L첁�j	u���=��O3^��}g�.��9a�E�EX"% }+���酏�Ci����|��v�1_þ����1l�
��ER�.H����>�;�m��u����c���`�>?���S;�I�������VLۀ���@v��"�+��y�溬us	�m:����`�0����{XGz�5Λ!�,%F�o��%�	��\C
;�%8��]��Z�6��������.u��_�}�2͞gF�ΛR@�u�f�?=��_Z�KJ��z�kӶ��*�N�Ғ ���Q��!5E�򌕼�%�:!��w�à#B�VR	�� ��w��&�5lu��T(&�v�6b�V�nm�Zl%$*���K�@��%����N2�$0�������E��\7�+�Ǝ��U�%q���gǣ�b��F�W_�:����w��v1'�Nw�Ù䍪�]�k!t�z`��lԆ�5�I,��XkB�N�,�b�>����@� �7��?U9����ժ�\l�k��hU�f�D����""�ޤ���K�,�͹5S��T����K.3}
~mm}"M� ,�qo��]�ߔ��2�l.��g���p7 ��u��2��ґ]�ڂ�D<}�G逅K�Y��c}�_�]��̢u��E�6�O�R�5�v��E��@ڢ�,٩���*c�bbŧ�Õj��rf(bF2�5�G�a߀4@2E�քK�����p������z���i!_���ܱ���W��2clù.�a33�@�%F�THZ��_u����l't��qfQ��1���PXa��ϳ֪������1�$�TBˢb#0T5u\X}��U�*K����gO�tgh(��K��+�y�ju�v�n
��`�α	Ȑ{�{W(�x��:�P/p14�Æ���R��"��%!K��c{�:l�ͯ�t�Q\��qك�y]�����tI����)qKI;��(u8v�I�S�Z�uR�md�t�۟���::�S�һ�ob��D&�{9?��C�kR5��5!a��v�N���ψ�CNͽc��t��P�M�CZ�E�#��Ô��QYM�Fϓ�Ւ�%wp#'���%0[e{l��g�/ds����`���Qh�	dF�G�Us]v�$��M`��$ʃх-`Qj�2�Y�_�l��	����C˃�z��G���^��7�񇢭��?ۘ
C�I$�;B$ �Iԛ�͢&s���ܱnn8�	�8�1�`�?�3�\<�ςx�qd�+-���C�.�C��%��z��f��F�<By���Y���$�UUYc(�2(�[�WV���x݇��	�
3�E��_ 0˶>3���:��=%J>��*gE�E(�&NA%D�K.��wVϳ�rJ��I`�Ȝg�����wykv)��TB�֋�M��d��������.JKв�=ݦ�+��6`T{c��l)Z��a�P^ ���ʸ���tx�0�׫����y}��CȥD��-�^���rRv��pj�������/C�%��⯘��4t^��Q:���)���r	G�ƿ�*`���C�+tKH�G���1]�I��G	�(d��]6&�@H�VB��:����7��	iT��G)*A"���4�S����JbB�j :�����\�v�f"����$46z,��+S�C��N���t�?�\�rm�<׽�t��� ��!�t� ����U'WF�S�a��û�����3(0���ƞ�J�,��t�'��J���4x	��Mll���W
�V!(�g�.�&N������2�ːY�$�>�����R�u�O��$�ͱ
β�����A@(�~s�:��V�Z�v���AS1��Tp�Rs|i�x�ڇm=Ϸ�z���g�z�_�	[��=��x����ͭ�Ww�A�b2�tSeMX��읢��_�6��4��y�����+>�̳V��Y��By��X��-ݝC��xztҴX�
�H�S�&���w�CS^p�׶��1������i����Q��C�E�� �����l:�,��G�q�n��]���tl�qf�
:D��Rޱ�f��o��R�KK�#b��1�;u����a<1BȔb�?.��C��k���ZWdz���Y�v8�Ҕ��F;���pH�bi�9aP�S۵;��o*���0×����_y��G8���:6�zp�^_L@�
צ�;Q������A���g�=̺������8]�y.ؽ�7�C;`��lp�*]�T�mS\���vO��s\t	�*�-�}4=�f킊�P�t��e�0�QKі7[��Š��v�q�}�d�d50JB/�s��I�������p�F��e�X�B"%��p��J�i��yi>���y��td�Re�)n(�|��Ӟ�X�j� ������>4���6�k��	g�hk���-=@eV�A��N��k�Q]�#Wk�O�q^�ڃK�]3��*YM���)��;�2�v��M�s��eo�}���EumLF��&Ҝ�8�	Xݼ$rHw��������s��j�6/L{�W�X.Q�f�ܯ������d
���ǉ��u](��"|��|~_����,J�Y	�Q��ڻ?b��fݫ��"�%x{��T-�l���O[��ͨ?���%^^�u�i�v �ъ��.&n�.Ե�S�B� e����D���ʸQ�D��ך�Z�b���"?J�ó>$%H��s5�hʫ(+�Z��A�d�����'b_��oH��T�ee~L�cM��o9e���D2�r�W��)�h]���������e���iv�F��sEd�~�u��_�C!�O��������;{-�0��*�K����@Ws}��#��S�;O�+q��貤���5
?�J?�����,��Pq�2�p��WFrե��es�C�O�22�� ���K��W�xg]W\=���Hs���R
5��/����e�ܵU�����m�B�<h�G,�>Y����sM�e-�}�֎]#���b>����J�p��w�����.nF�."��P7+t�{�Of-�ׅ6tr���K�QZ-�pO�x�8��3q	폩�!�����_� �)W����m���'�鵛�|��'�{s,�x�;bN��YTy�c��2 ��V�5]���Rp���p2��0����nѭS8�Y�M"��"���W����"�J��^'XlT_$��l�Z���C�,5[���F,uzL�6���W#��碜65��[g��{ }j��Ob$:7LG�?�1 j}v7y2͑w�n��N���4{l` �66�s�����I�W�Z�(JHoκ:�a;Ůd;!�sT�
�I��6lP�m@��-��
����V�	�#М�}��˗�D��.Ɛ09�5�,�U��CW����
��?$/$�������	_!$�-�/{bfe%����ǉ�~d���R�H�=օp�!�07�Q�i{�X� `�%"���x=�zb�>,�d����A�6�&�m����Z)I��GAO��+��mfO�J'mθm�p��eW�c��+��g�]��D��)P��Q��՗�X25ń�*淭qmv|�����"�\��Z��z�D�5���	���Q��g�ޅ�p�x����L���=
xe� OQ�c�Q1I���*;�"I�	�13C=�z)J��<�w%��J,�݀l�{�fdT����|:�ۑy��Z_ʟ�6��ຨ̵��))5� u
��q9l�"����	��yv�
 �s�"�-n���^���)qQ�;������2���kY|#�Ŝ�$�M�i���7�VC��?3����5?�v��U��3�%��T���:5X�3b##qQ<(��e�%3��
��#E!��	 �\:� EC���'N�{��A��q��<b!��/��ڙ�ޮ�0ɇ�I����v h.Yj� �A��yJD�r�i�4>Fڝ
�I\�P�{�3t��މI���QC�`pb�)禃��AeS���M�������G��iW�0�g9+c)	�R7�L�;?#�X������F���X��I���j~d��ێ�+	L���+k�/��>=θ2� �Wt���3ɏv��T0��t�A^Ց���&hrB_��X���=��)��3�Y�>ʱ&��Bb�#�W�������A�"&������t�	�.A}���ӆ�K
�}�v��"N�*�5O��!��,����>ՓR��r���F-h���LIM3�N��E��逹Hю�7���������F�[[(t�~��� �Y�5F~�1�L���ACiS��E�s��l1B>�W��zR�jl����JU�"	!��u�&�	ahl�k����\?�.U{{y�7OշMA�1~\�q��qL^?_[:��+���=S�9��f"�g�	�JCTFłMՕ8��������:��I�AI7�©�T?>JBpހ�.+��tL4��6m�r^4^�$V�5��$�<%�-�F�1��|3�2TP�@>���d��'�v�N!��~D\����s�rN���E�/d����p�f���tݥ=2�$bS71��?�f�W���ߞ�>u��0ΐ���~n�䡳:zT�k�����8�f����﵉�A�?6l��l}n�?�:U5`V�T�n��ǾE��9;R'X�L�gnnF9�%�d��^�qb�2�d�`�XZ��nVI�?�z)��+5�m�s1��\ V�Vd�ݐi�?�f�`J��L��en^��g6+�U�:36��%�_�p�H5�W��̝��p(�;��i��M��Ӓ�\}�}[�5�{ܰ3��.��e#fi�F�J3K	����IO����#��+1�5��ݚFl�������x���oH�J_js��b���4GoQ�<,���@��r����9<��p�`L�B�#KF�G)����<@u���`����������ǡ	��{|a�?�j�yγ���T����Z�=��j��J����²R�+�k��]l/CJ�Y! � 5kf{�|�5|��g:��Q��	�m�3 ���s;g�E�Z���~>�xqS�OB�i���z�2e!n�^P@1A��o�Da>D�Z��g@��d��r�@&�~$��R�e��.L�Z-�'�oj����+���ˋ/=�kԐ���s�9	<5s�W���Ԏ�7�/k�s��H�%
}TI�f�i8��T�5G���љ[�=�̜����?=�6�M A�h����丸����V6�;��8���qUN#L�	�_���ZD+9;0V#P	�P�im>z#?!�Y�J�0��Ϣ�YC�	T�4ъ�b���4��8fN^�Cw����d$]���SF��Y\B���n���I������**�$�~mSJ�d�8��'���?�r�Edd>�vS]|��կ�~V���h�&����,�K��Y8x7ׅ��'��K@g6�w��~�ز�@��q���8�
���#�b4R#}\*���ٴjd��P;�I.��|�:��1��p����8�����	>�das�B.���e��{�?�A�{?=��Sx_��.K\M��|=���N���5�B�b�:�[d�V�أ?p��Y PЦ�t���_}B��u� d��_��T �Oi�lR�������גx�)"�D����`�h�!�o�7R�[E?z��V����V6g�n泂�M��a�����8�nB��2T��ƿ�z��oӞz�P�c��Z���^�j�	����/w�Nz�3����ſm���0�M����^�D�Ɏ��;U�#̤+�Rޢ/}�;�L��#G�P���O �r�.C2���P�{�%敫tz����S�\�0vL\��%H�AB�iZ�8ض� ���2�z@��Xz�?'���Eu��G�69h+}j����-��KMe�$����	�}�{bJ嘢نJ6Ԃ�I�E�δ#I����l\}�+�U�/W�  �,��˧}Q:� ����`�Š��u�vW��ۭ���W/�~�]��?Ev�_��vvZZo#��|3�u�d6%���7H��~ ٘���\~<��V�1��Ɩ3��;mG�������Iǎ(O��RV+Z1vOb�T�8�h�a�7��KbkP�O������|d�"m��!} "����ɞ'?7�*��~�WA��IK9#���"ڴ�Z��ɮ���$��7DL]�Z��AP9�m��o�>[|-���m�ph���{�.�W-%�Pt����z-����)�wT������;p= ��
Ī6x�ը����3{2�'�49��-1���y����9�mb�qu<_�]�"�QE�Hj}WKw��5j�W��c|&�C���}�2L���o�p�\��O��1g��b����l�M�Tn�T6���Av?$����K]��e�S�����ZZ�_��� k@���8���ۢ�z�z]��w��5M,I�B�t��D�2e���,'�}[NMƴ��1�bG��r�!� �u�)��c�Kx��s�]�f�8K�����Tn�9�aF�(S`��$�u;
�F���S��c,=��G���b^U ����%IP�@K��1M'-��[��1F�B�!��ل���$l v�C�j�A����`~�Ľ���?��� ��>U�:�3,�W1�����D0c�a��L�]\��ɂ{�UAvhS�������ʀ�y'G�-G�)*"b*�q�
��'�C)x�dw�T�D�pwP3L(y�܈"�M�
�KL}�4�YxCfF�b��@�2�9�ρ�؟4������-����H"a�Wn9~f�@�Q�Ւ�A��-{��AS�-+���^�$>7���Gc�=o%kLIhf����xX	��9ԥD:m,9*0����&��x��J�X���4	t��Q;�'~$g���g�"�0�#"�}XO�$�|	�sD���d��`��F���� =�o
'�������I&��e��6s��N�Q7���Z�N9A����B��8�[&�%}��X�Ҿ��Y�B��CW1�r�|�ٚ�&��R0Vq��>
|	n��p�剎�3�]��2�@;�ϦkmT�HOh����O�IA����"�?���h���g?��NV�sŵ,Trv+Ͻ�
&��j)D�h��"+�k��7G]�b�$x�]��;�7������:�+9�6��B#���8ˉe�������2��k�+�hU�8�9[Z�L��͟"��C S!�%�j����6�%F$�;�s�$r�呍	��TJ�Z���@>�αL�i��Hԟ�p��϶| ��l�JUY�'�:U�3iXrVK�|(~G��pQOw-f%b�}��D��M4P@�#�;��!{g��4(Q��4���YEݨA��`n�������|R�d&S`��8���m��>��<V�8&t���j��7·$5�(t�������N��v�xH����u�'o�A�y�3RJAy��& �a�a��[��.{!?��P�޻�%��_i�2��t�ݷib}(�����4�>J�T�6�f�q)u鐃�a��%�!��QQ����������X�?r�Il_���q�D��x�]fO9����@D��������l�Г�uI�(�3�D�tS]��j|TH`Ve�M��t�P�:f�����3kr�hP�;_%Fv�̅0�|�E눇�`Tb����T*�� ��K{n�e�,����6Ӟ"���~ʬIP����;��TPO��U���7d�����*_J���"��zp,#"����ށ3e��K��`�{挗�T�c�S��X��/�������}��3��0��TÕd�f�L^��j��@���p��|���y����{o�qą��/�.�	���:�"/gtx�R����P�H�e��X��� ���3��O@Rb�+�C�l�R�����ذ�"կ��e	��K
����5�����V����������1� �c��"����#��x�'W���H��x������
u��[�$%|:ؒ0�\�'͵��p�EHb����ح������HV�O��YCΣ`������ا� ����F�ّV���������_����9�d�"��b��3`��		���=�~�UKl�����|��~|sx�s���?�P�F�n���{J��4�NU1���r���[(b�3#���c� �Wj���%��`Yoi����Ǭ��;"a;� nBD�y���+&��Rl�N3$�X�Q>�G=s��W,��"�����-�Փ%��D?��%&�W��j�_{��
\u^�P���ޓh�"K'��t�ȥࠎ-*�:%(|e�N�r�-J���Og
������l�Jx��@���r�݀�n �^Zڠ�� �uFB�9xުIr��R��!�;��nս�'�s����-�{�,�D6�J�:ɹ���R
,�>١R�gb;���M�ѽ��x�2���,�#�JoN7�8
J��D;Ⴝ;��졩|jk�&�^�[�̢� ����i������h~2!\�a`ZDE�����ϙ������Sm�z�c��^��іI֋��F��/b�r.4w$]h{�Z���&/��w��y4R�M8"Y���7Ă4)%�����������Ɵ�W�@<&w����wXQZ5a�i��[�D��D34�m�V<�N�6�˺(��ȶh����0�RV�� C��SX�Ĭ4��u7�[�U!q��M+��/-S�BL�1�Q�0I�P��.w9sy&�|��E+lg�ܹD�lR���
��7O(1ED�I�/t�:�#�)3�Oz�f�?bӽ�<���Pψ�b�<���ꚨ�k6�n@|
ƕ�*�Z�<I+#M�'�+P�'�D/����p*�R��/�dD�/�Nѧ�[�+��'gRB7AE�>��-��?f�a�����c.E8�֡�٢��J�u�!��C:9�]jX˴lF��Y�|#lhVhӤPd��Z�xp�y/���	�ڧ�h�m�|�s����>�駜�$_I�~�9|Tm����
�`�ټ�1Ew��q���Gx�hm.ڞ`7���TS��c�n�ɥÏq�Dq�%�i �Q�tt�T?�)_���T�]�}V�SSC@x[9�z%L&�1�u߫I>�$^�X*���$34���
�+����Ӊ"V����?��:�%���)'��x���C}�rC��Q��
e.L�����֍H z2�����,�0J��`Q�,�x�m4TKL)��Xwpm����M\��뉽����P����&��8�p!I������
*��V݌W���\-zf�����ǜg��~�T+��]��e�O(�C��,6��S�Z�y�*�nz ��:�?���G��6r~�5�������LQ����ҁL��"9O�j�h�{�6|r�'-&��?f�M�$B�垮y�i&w:��"��Q��i�9��VG����&f�������_�9��l�|�&he���V	��dɈ�)[C�<��lg.��Y���J,E4C�� s����g�c@k��yN�Pm���T�@l���Yb��U�S7@���l_��s:Jw:�M��̦k������3�I�/)��n���%���Ǧ뇺k�vX�k��v�u�MHf��gJ��g�e�����
Ɩe�j����L ��v�i::S�K�W�4X8���|�]O��B��U�
Aݗn�/%�F~����SH�E� ���� ������I?
�ػ���{i["��t	,��8�yo��v�j���	�(n�蚼�j��oĜE"k�g����W>3���^�Bx���c�/�k����J�N	(J{c��q'ܷ]�S�71�Px�nj�}���j�o����/'mQŹ�&�p��sڬ���(|ɪ5+LX�-#)e��x��{\��%�L�H�Vm����Q��j�2�MbLR`�Joh����t3*2�T-u�"HW:Z3�٦7y*�[F���L�2��.J�n��Kv��B���N�T��F)��P�V�Mш&���8�1΢�\�u���q��H��v�c�ԓ�8d�e�f�ܜB�7	>Pd+�g$J���ׅ���i�)��i�.Q��>�ʹ�Ҁ����7�sF�@��^n�'B��djDzt|Ă��t����'��=��/�/U&�Li����/��iu~oFd9����!FORU<+���r�s�9�����+w�2I�0V��4,�������r���IȺ(�����h�*����y��b!�� ���%E��-�SqڈrDl`�R���TT$��l�>��N�݊�Ԟ�C�ͽ�j$�q��Cjq��e̊t�Ҋ���OC�]�E��u�Ks���j�uN�#�Y��"�K�ꍑ�����*��Wj).U�w��rQ��-�D��|�+��*u�{vuI�ڔ������K� ����m�_���+,����qSЃh�3C��l��s/�������>���+��N�"�:Z�lP��Xm* o+��e����­���3m��N�i�8@D|�2�R|�#��l4C��p@X��]0z�c�^D����/,�zo8k����^��$�z�2��C�u��}�b"�l_*Zn�QU���R��)���s�$ ����=��/��[�vd�QxG�R���+wb�%Ɯ�pJ�Y�AA���4aY�ҬM@B��3Ɩ�[�ڨ>,lva2<O���DFH����g���g,�Ͷ�N������<g�,˨��܉�ɿg8�vq�?�g5@��=�@��1أ�Ǧ��_p���O��r��g�'�5�a;<������m�A;	N^O�i���hUru?š���W��.���]z0X?8��pkF�W�D��'�7�~�9��+�f�у�!������BH���߽7�iZ;�m�:�n]88F,х��E`0 ��+r�zn�NYeʗ&�&S�M���W�_�Z3k1*��\	��S�O֗�,�b(:�A������/1��;����P��Ei�<Ȋ{LG��"v��ϒ�M�ryT��O�a$OB�)H�5t]�a�Zu�����;�� ������	L�d��~��C��5� �<���r{��W��N��u|q�!�[���(�x;����&�AἋ�����z�Q���^���m���P��KU}܋��:G�D(�<^�?�|1���Yu�L���4��8� �`[.좌4�^���9��_pV�&�)�PD�X:J��*}|1�=)��Lbz�5y��kX�C��2���lX�w���U�w���dqC�*|9եR;u��)�Ci�d�d��x�K ~0Ս�N����@5��n���j�GS�8m/�N�&@cjs�k@�&����
ء�3��j�� ����� (�p����<x_9az��3�y��T7c��bݩ�T�ߨV>D'MD�Ҽ�����#�rr&�����Xx��|d7/8D���jҙV+�7G�̢%Ч�ي,��@9��uO��Dڱ�Je��zW �Q@?��0��e�*ӍgE4���������,L�N�h�^��͛C��A{� ��|^�G��n��3tʥo(�l�a$f�h=��!�rĐ)��%�x׸����1�< �"��ߢ�� ��)X	e�����?�ֳ9�R���G{W�R9��1��Z`�Mx���?�J}����I��Fn�Ü���vO~���g54�@FsO8.�xOF��+�-T���m1I���%D+�����IL3=��l�mE"Y���0v4[������P�7�M�-�:��փVN����S��B.��ոR��$�8
ľ��6���<9���ݵ���P�ȕ���$��&v>��%a?75�v���2b�@��H��K�a{upB��Zwa8�l�Ɉ@]B�]��qģ�F��dB���?�*׼���	��l��G�| Mx�}ֽnoo>�w"m)|��t��J���gmG���o���1��d�\�(&MPV�~B�����(�T���M}��;L�i`�ܰ�2�o#���4Vw�,�BH��!0q	=��t��kŭX`���ʾ92?�45Xٻ�ތ��Cy�\H���fUњ�����f�Y��\�""B+��J ��ӆ�8�Ʒ���2ŕ��"�6-QY��,���3�SLT\7 �?M�>�?��0j�$�:�\�ϵ�J�`��V}�7%����qI�8Z򸾦:���;��T�:$c;j#�QF��e`۱�f�d�5��6@ �F��^k�'�pc`�;�$����u9��2���f,�6-�܁a�$o�W��\�����pS���spn.A��|�i�"C%^�K�ʻ-"�H�~7�x��w'�Zj�d�<Bm�3%r��n]����}qs�+�l���FM`�u$ᨄ!��{D��;� ^&�i�����0����խFRw��| �A^�]���Vm�L	9�,�b�����Kb������%c�Q����(�O��-ekD��3%�Y�[�c��Z��%FJ0A�m1ڧ�̚�٨N����f������C�)T�y�ǃ֘���&o@?)q�ەq���[�}��f?=��0�z)F�����Z����.;���ZWL��FR��B-�z����	z��JWw��ן����	��nS�J����/P�	��l�	
I���Gݳ��=��Ր�O��N�h��>o���xG x/��#�e�ڇxͶ;���}��v��0���,of��p�9�R�r����zة[>u�e�oI���s�;�y�g�C�O�3�P!�����u".��������ԡ��e~洫�!�f��rQK,�S������ZZ��n\@� S���R�:t�na~���˿�{��	�ϰ���3�w�τ&���]�f��<���T� ���^�t��}PU��U�����I#�M��Ա	�Lf�H*��$� ^�8�c�m��Q��|S�P����V�7���V9hJ\6�.y�d+��%��� ��>M��,�6R|0�E��9��i��(�[s^ǛًPy�*�+M{n��[���&��g���J���ws���q�!��8��ls\&/;\��=�ou��s��|%��B�K&�-��ƈ����FՔ0-f��8��g��UXM���تai7��a�|�1ikm��	���n} ��ti�����Yj��xf��� +\Bt�����Q@8z�1ʸҸ�ݢ�n�pQ�N��i$!�  x��7���v������tUl�3^���jE@dr�	��+�w�O���c������h��{�wm��즗�q�;�R#.ɣ����%��dל X�~YAK�Gr�]w"�+Tj���^�g���W�=ό���×o�����Fyx���g�>R�âH��2�m�*_�aG=�/t��S����-x��{�f2�VlXTTh��i�vK;�� WF�*��x���/�$�O�ju~�#t0/�~d�`�O�0��Vǁ°�K�+��'X��eAWFv'��\�H�MM`b��th��l<>�dI�r��O��+�zJ��5o;��7�Wg������ǒ<�m�/�����y>~UdX�?��f�ǩxF�\*zo��&���T.�
�]�d���	�O�rۺl�K�������wfh�	�]�ϣ$��xM�)6l')��ڻ�S�����@�#�<�\}�I�ʛW�zhޡ�.kGS%N�A;�F��s� ����KYbs@c�V|T�ش"ȟ�酌�5���M���+�nD���*��pOso	Ɖ�;$i�I�d�l9[Q�C,�k΃��	��7���SB��!�/��mi{<jjA�R�`��"��[�������|L�K�_���A�!Y��lGfs��˴ޱcc!����1��O��	dN��Y&x6*!Z�]���)�r�Rh2�F#wm�x���ء�]J�u���ʹ#��VMw��gu(D�*{��_�R�8�fւL6���{��0���2iGd��L����?��c+C�t��$��4,O(-kdfpj�gP��6���B{2U����=

��i:�����w�i��_Qa`<x������2nR_��{�5��8^�t��K���mgU�;�$n2�\����|i�X`�����L��YE(>�$�̌H��"&&���N|7����~<:�[A�/��X4�J�ֆ�%(����{@o�W�����N ���AՂf_7�	4��8a�Ȁ��xb�#8�!��n��@���+>.>�ި�h�7S�yb�̌}I�q.�@흶>W���K?�Z�Y��F�_�DSA۲���xV�l�5�� *.a����ҧ���(��C:��v����̹ <��1�Y8��+���ߪ�ژtj�~S]p�PЕ��ѥ\c8p:��/,J��=��Wj�ׂ�v����\�u���aҢI1ڬ9�)�~�4új�ʱ7�1$Z7�b" ��!+�I~5=pPq���������`9ѡ��9St�f��s�0ɕ@�س�c*.�uҥ��P�+��8�m�Ҷ:��y��l��U�q� �0�H�X���c��ff �SQ�b��)�v��(�����T��V�Url�{s��Q�7��^SU������#O�����h.�+$�%�:���C��[�u�8�ș#�ݻ!޹�7��q�_@��9�i���~�ٔx�m�.,��ַ��.�ݡ8Vg�]��ʥ��k����6-��0�z?�i���͊Bnj���
��[N"3�!U�.�ś��nޙ���ퟧ��7�}	��W��0��܅
�6�קu�l��^N�#��pQ�pp��
T`T��ɕC���o��՟��4#b]�BN8#�v�(��F�ۢ|k���E��cyU�Fk����_gL%�fϑNM�7t���2�u�Z��z�*��1��_e�#�p��Z��1�J`e8,C�A��V�`���ug8įj��n��؆�L�
=������B�8�D��N�p|�����C����;��~13�+�T
���??)�.�{kʑ��̡K�/6�M��y$|'
�!.V�ܔ�fΘ������[cv�,qQ^���g�Q�o���JL����������������:U�� 35�i�p��rG��a�{������b�$}K��.���z���H-ds�)�[��%鹿%W`��S�V��FңVUn���+aĄ�xH�~�e���J�g�
�E�*[���m #56����Rv���!�<簼�2j�b��+�Lio?�d�'D{�	Je GV���x!�tB��'r��$�9�k��]*�Pl�ۋ$w���뷡������B|w}R&��O�J!v�e�u��Jf/i�(���1�\^�+��^R[Le��KU�Zʛ{��bS���a_�/S��Z��k��y��z�;�k�tm��d�L��+�e�J��ʛ����
�H��N�;P���#Ư!��?eKԓ�{��	z �����Ee�ϓ閪3�)�e��VZf��C��[�Y��}	j��Q��?z4w���aVM�[1:l�B�`�`$;&�Cщ����
U�p<���9cƜ+�_W)2Lj��j�.#���_{/� �@�J!�T>Ey�8w�?�V������<Ж8���i��,�g���_�rW�)�1¹&-h/�����'��\|I鏴l����ϴ�0=��p��MaB'� ���!��
��#U�<|3��\"�;x4��_��x�^;����eJ��t�Tdt8����W=FVp���F_l�'8c��h�7����!��!�6�P��~u��F��y�m���p0��M�P��!�D�X����`Gr�%p�԰��%vߘ�3�}TG�n{Pܿ�^�hj���,�jךּj���0Г���;�j��,B�ds�vh�D�g�S%��U*�
�����X���6u�g/c����Wi��b(��<��؆9W�Ʉ�f*+>7H��c���{$��#:�l"��o��N�:c������!�z��	�se���g��;O�����x���A��4�Mr>�B
n �uj6k,q��2���M���`h����Q�78m�w�r�Eu�S%�@@�0�1����2� Qj��~�Vz�e��o~YֵٙW�.�����#	" ���D *�U����)����m.{ݩ��_,��ݸ�\��_�{_.�:�*�N�7u�/JG���aJ=Y��TНt�Uh䀹d�3�k71
����*�Hi�)-�z{U.��#�׵ b�)��|�C�u-�;�X�f���2�h�W�=����A���@�^�\t�=�r's��6V�ba[Q!�+#�ޯB��� �����.�W
j���9�9���E�N	TP0���w�7�f纍EDՎZ�po+�%����Y�L���� �^phjK�t.�I�ܭ{I�W6ʎ����Q��dn �)r�����k�q��8�Y��	�6��M���H=�L`�÷#^:��`Җ�?z���0 4)�zh3 ���l�B��m��M=%_�M��v�
��K����m�ɤ~i��Y�x��r��i�r�*4��M�a��L������pD�&�s��z��[뉊;W�8�zP�������|AF�y�G���Bv�֓r���[�$k�vD��=G`�@��G)9�aU)��$<���O���hUn�C4mQ�<���䑺�-*P�/&˘j尅��+Q���n��ܨ����� �D��T�}E\��|�ɮ5]N�֮6�<�t��T�Fmd�A���mj���f<1=��Ydl��kz�M~s/5$D�$�Z|�l��$}����ˑe^�����u2�� 9ť��H"�I�1-6 @�X�����zD�[��z�9j7�?s5V�U�B�l3��WuN?|4�m0�L�pR�ip��H����f��ތ����bf7�����<��7S �ȱu5��=6�e����HGȰ�
3o�N� ��VY�G�uL�A^&D���bA`=~7}�]4ۢ�FHo_kd瑣'n�7�K9F�lQG���ΓvCxS��-��m@�2�=�̡"�UX�t$p3�̋ �3�'&�A2Z�}�*�nމ�V�J3rQ��Lݯ������c���5�Ȯ�QQ>��Os�%zTj�<M��$޸�`ڽ�zl<��3va�����u�<���C����_uA�p"�O�(K�/(=ri��b���]Q޵�_&1��B�;� 2 ����>߁n��i�c�Rpe}�
�Z��׉)���r��ZzD���	m��ÁV�k�;�ւm���z�?�6e�/�J6���};b��I[����묯Cc1	����-���4r��ڭ�ȡ��ΰ�!JS3����h&��+�_{��u�;���'CaJ�)V[oTS�V6���nѣ�i��5{)A?,���d�$��0���)D"��
��}��� V�XƏ���.�I�_�RΌ�j�+�rB;�b>e�]#Pf��-�L��/����kd�n�[T��F�&��O�����x��b"���\��Ts���.33/�7���U�	~����%�nDڐsk���^�]��
m���8Q+@�A�mm�J˓�A�V�݀t�� ��d������w����`�_���͓�7t�X��,eͥ����j }��t_�F��Է��$3E�ZQ�{Yu�*'���5G��|1��cJ�\���&HV��Z��`�ݫ�H�L��Nkl�7���)�o��J!�`Sb��?X�bլ�~I+n��bB�M� �l��s��H9�-~��v9�}U�۫ST���W�tV�0Et���h*s��يx=E�q��5�Ȝ�����Dp��-˴Xl�?u��x��Ye�;�V.�{�l�p�6$ZeTlZ�%a(�d���}r�W��X�)�����2_p%8�Q-��ۤ�jx��&+e�����f~aLTbh�?��� �������zZ���C�!��]/��[����U���ڒBOĒ�,�[Nv�����N���m��U(�M}+r��i��@�F��L#�<���BQC�� &y� )��x�m�@a��p��v2�9
�F�j��l�D7�mw�i_��u��͸v�ű])k�t?���-� �O1&n(��[Wc�bzӈ-�}�s;�$]��ԣ&��/�	X�!��x/?���knmu�Y�xx��v�2`q5���n��#�泷G0��(mS�4xUyx}�{?����H)n ����qCV�А�Q�9<�ۻ<fl�?17�����p�u���Ё���xn��"�>v�2�
!�%�v#���1�B)56�?�*�G�(W�!�𸦏���M���-�{i����M��
��Ǖ0wÌ0�DD������g�ƾ�|���~�`Å�A�"��i��5N�����5U�aq���D�^�_�T�6�>��{k�QL��������'�Su�!:}35b�:�7����;*�4��5�n�{�6���e�\ ��. �$�`�g7��.�(0R���]aB������h@����.�9��4�-D4FBQ#n�ӭ�Tۏ���e�r��*H�f���Y9����V�� B����rPx��R��IQU�ں<	{��_M˿�3`�-S�l!��s���Fy��(#/eV�������ON�H���@n���[W�{ B�r�C?Ax��^�����ش�'Φ��zSj�5|3H�\��0�����5,\v�!t�k��tY��"w�+�u2ΚfW��������E�,p�򮞄*�?��9� �#���sD���R����݅n�,r2�����X'���|杧���R��=#����G.�bKW�F����� ��d�ӡ(�¡���Y�_z;Y�U��/��RL�5EW�C�h���ӌ��y�ur��
��*2�\tYU�D-���;�W�LaYvt�N�Ŧ���NU"�A��u>m�Z\�WCY�q�U$�ZgP��8���!��&�i@���r���\r
a}0L���߀@����?�{���%�m�B������vŻ�#.����Z���6�8W�մ]Q��貝�5����NY� �(�����H�����S��XԒ6	��`��2v7�b	,rˢ��&H�L������������F�^�eo��ϽƱ���D��FeC�����'�k3#�A�%,��Sܿ��Q:���_$;�j���;����^1��t*�$�+� v��5��85��gLA��HV�S�˸�6
4�*��E�\�t��؏hCۑ�]n4Yk��<�!~�²��/��H#d�q��_J���U�F�/"俰c(b���o���SR��Y� �lR}�<��N(��J������Dv�Lq�7���[�i��#��H
Bs���Ta�|��C,���걤��
$�j���BK�ziJY���y�T�\�9�i�vī��9�=� �qo�6s3u�"��G��m�T�<Jx��4�@��!�}��j�y�xM�A��9����	+���� �d�/*+��/#[֩��{�$�!�8��	A�_������'��?�m�N~�f�vf����`�<Z�����K��5_Z�W�Y�Tʂ�r�7C8��h@��L�fX�����Ae��F�9���ZzI�pv��X I��Y����2�8�M�4w\�e�_+�~�@�%��'LX].���C<zC�	p~vg�~��.9����&�d4�����y��84gV��=�0l1����Ț�,�tH6C�]qX�>�Y�%�#�S���o|exHL�QS:�V;�j�����0|w�2
�{�i�����x�@��N�n���䱼!�U��,���T|d<$l �g��\�5u��4z��soC��0�� �hluc3a� �L��{���,�T,|!��ߌYu�f�	�PS%�����i�r���oTrQ/OK�\���	ne^�Ap�<��Ш��0��2s	����=W1�'��X��Z"\M5.X�����.�1��b�|���@�^r{�I4��$�������TV!辫:#�,l:,���V��G~��m]U�X��� �$�Q^GDz��y)9���*��q,���
�,�����XR��C!! �wZ��"�@�'��S"#?M�1ǡ� l�X���Y
s�(�7D�S�.��$<bv�"�6�XQ�:y�s�YA�� ��u���n0��g"�K���Q������<��C�Ke^<һ�[�n���\F/��?��z��p��xyf,���]KS�o��\�J�_�~�s�V���)Uj��}0h_��>Y��wYd��3��J�wL��Z�C�6Bx��5 ���}���u<z)ʫrr6����t�F�2���<�B���w-7�1|��B���&*{q��[[��p룯]�w1@s*z<��Gz:���_��c~	:��9|������5&�^��Ҹs�d�r)u�q�Qr�'�nʍ��}��iI�``|i�L�h�KIj���dL�r���x�/��M�T	.����	�;,R���D�-�`E�����p�`�?ȠQW�{
?��$p�BCڅ�Ϸ�V�ziȲ�E��[c5�9�+�<��ɋ���z�� f@
��|]����"&�Vu�1,�����'/�����N��l��0�BzmX0�pd�8���ĬW�X�*�u�	�;j|$��6�^��hoI!����ʞ�c�Z�3�%���R�Q2�ݼ7ի<���3q߬��������u�&u��ܔ�t����fW�g(��Аb��	Q P�0Olݚ�58I����"��VC�n���[�j�ʤ!Cћ�i�1�g#.>@6N�����+�ѹ�/�I���̻�ԿR;p�U?�z�n"��veǃA�!�q'"�W�c�*&�!��N���/t�)՘f���d|r����ө�n0/XYZ$?l�;�#����)xR�k43�_b�y�S��U���
��x<�t�H�N��@K��^hE���0!�0./�֯�H�m��b�����3�<��.*�ش;y؈��3��o���¡5-�ئ4��/ȩ������r֖� aH��9���U����:y��4���g�� �$߷{e�?��Y��~9������rH^�!S��4΀!���U�W�"l�=�T���MV����q������]���(-��pF�_��vnO�P��$���*�C��8��u�*�B�m�
�����s�/��8}������P�ܝ�<���d���?[�8r#q�����u5��x��F�)�O����Eg��fD�ү������_7��S쯗����(ҽ�kX�[>�f��W(�z`L�Z�HU�P:�¬O+%z��b�N5�~��١̯�G�:E���9C�V�" �<B�W�3[h�������������^}���4�8����>o����/���.=���y��j�1�9�o7���T�`q�k'b}�j�b3ŀq v�p������'��Yd�]@��gT<�����}�l���W$ɑL����>���ki�;:�K(�]N˔NU�����GO�4cU�_�(�������+wP��^/�WEWcL��CQqv9�(�t>=��?0w��G:�F��W)9�Q _OX5d&s,<����Y	���x����R�"�`��I�~�7��eB���C
|:iF��,���7wT31w���.����R���P�AuӀ\6m���G�g��M�|z�b2��bAօ��Ew�Z��Q�txv�$�}j��ߘ"Ȯ���
F-`��X�/�0��	�F:��
1��\y�Z��+�b%��fl\���jiNOF��y�Y[���&��WO�R���' s�<�qy�Z~YSJ�Rb?��H��?Uɻ��G^�(_hmp��x;;�\���|�q�jx�2�?�V«���wJ9d�h��^��J�Sn	%\`��0���|G)�ħ����O�9���I@s��_��Y>h� �-�¼���f�<>i��{�A��7�Jn1,=�r��LU �Nu��G-}m��B��O�+f]�D���+�j�I����Wc�����^4����ި���S��RJ����Tʉ~��r�ٕ*�a�%���lh��2Z�q�d\���1�X�6FÛ�M�ǽ#��,�@�w�>��BaJѿ��#%����ʠ��~���ʜ��.���}�&�T}�]���А���A�g��`���XN�P㺻*߁�Iɢ8���і�l�oĚ����N`c\��R���#\���cW�d��SGrR�'�Jz�5��g15]�g�������Ev�1!:��1%��]t�!`e7�x�n���*��ۤNM(��c�`9*�Mg*�R&�a�=�������~���*�	��,F�<�3rޕ�Å,�[e޸�&�������v;�]'�D��!�<����[�22�h���&X>z�[��奋Rc�hL�a�\/����%�e�=�%@faFјȻ� �X����ڐH���$�}_>��ӊ�#�e���{���6�S-55=ds-V�[���D�(A�+�@�2ǫ�=�O]B�B��Đ�2�гk��Ę��sQ�^PT��q�JIW��'�^%����._��tEb&"I=Rfɬ�y�_��ݟ�rT�k`)�S2ڴ����>�䁸������F�zޣ]L�8i7����M"l.�]��S �����l���P|~��o);�����4<z�NzS[JID9;�o�;a��Fm���W_��PIߗ"��5��A��&E?��M��]�� �m����9RE�}vX��p�R��-������r~���%�KT�Ŗ�v�gT�'Tq�e���&l�F�Q����?đ����U%*q���x��9X�	َ/�ʲ��ІX1V��fQt.��(,�Ec�b,S@.6Bj�`}�n�\��M���g����,ƵwƆ�3�<
��[z�����|Q&���/�#�3�A�èqn���3�.����r),]^o�I�2������#,���K05���U���=g�LJaE�8\>���F��g(B� S��mB�����Ժ�6,A��|h����=�<&��������1�ɝ��ڏ�
� �hd�pe�Q�HIn8�Qs��\�^����%���ʕ׻�� ��)�ly���)��h��5��x� ��r��0�A�La��q�-�U���cen�Q_a�d�;d'-#��e���Ql�������6s�w����[	U0?���Y:�Q����k������aH{%D�%i���A���3 VܦH&y���'O��LX����v^A�
�$�倓�e��Ze�A-m���`�N��h��]����Օ6�x�;�q�1<|�������"T���@/�}{�0��h���ا%�VΈ�4��I����\����9+m
���cL�l��yH�h��k}���-�*���M�VP��Adʩ�C!9�e2 ������ż=�J	��y� ����9�<
�*��up��82�yE����T�'��E;E�w��������"|�\#�@^`=%�1���$q�p� |�Ad���h��-+�/u�Qx*y��%�� \G%0e�`��J6`l�����-��RP�UH�:�L�*n�>Z�����q�.}� pͅ����DDz-�)6����L:%1�g��5w�AE(�+6Y��:n�[��f���+i��?�H+�_��X(7/�0^����ٟ�VN��!g�-��8Ϗ[N��/���0!�KOx���"���X�1͎k
��׵ o�
�N�bB�t�m���.�p�rw�9=#�<%���-�l^�(���?i;g����*3����29T(�G����[C�u�Ѹ�Ա�'����J��u�=�E��ظY��W�)�#�����z*dgi@gG)��36�0Y� 9�Au�dF�6j�s�i�Z�S�X?D�o.���������K>sF�D4Y� ��--f��.s��a�y�1���矸���}Z7��z/�QaX�|�JZ�&�L'mg/��c�1<�~�16�`^Y�x�h��^E�Ĉ����Y^��OB\u龅G�P�*���b���6`3"B��U��L�nPc_�+hѭ%�	��	j��bY'��xx7��jH�r��|�Wv�U�=�S���(�[W(܁y�'��zVA�����r@�0��@ݮSRW�!�z[补2>��CD����гhn���pM��Qi�@�n�]Z:���-��W����'�7N]��.��;K�U�N���Ƒ�i��Kw��4 ����� ~��n�{����P�"��P���Ѫ��氙�OQN3�ǹF��ʎ��a�y�GPm����h(�g�"�X%��Ѫɽ,��G��1����8�8���1�����`N/��$���zJ��i7-�@�R���H^~��\;��z[��ݍ��T����m��-�l�[���zY/�Dx
ꗦ�9A���K7�IgJ����z���
����@(N�Ԏ#T��A'��O�\�I#��[KO��Nrc�W���ʕ�����oj��D�5�lg���f~#D�Bq��Ou�>ƺ��
+C�Xf��n���G�߉EZ��߸�і`�@ԫ2�����:�}�ڨ~�X�/����T9$��� ༟����Ǝ	�IQ6�����
���3���ğD#Rt�����b���]Oe��52�ڍ`��o��x��m�]�
�b4�?��8%��J�A�ۍ�Oi<�Z�on�³�}+7G��~�N�C��X�,�m�U�Ȃ�*�u��Q?-=�s+K���(�� ��q�S]u2Sȯ5l|�t��=A�q�^d�4)�����
�17��%��$+��@_�<x�|�w����
�Y�LBe�mr��dx� ּ.W�3S��N^�$"Y��Ѿ��S]����j�hu�a]�R����L��|py��_n+�E�n���e�<
�"C_��9-�M�+!$3b���_��N�A����4���;"���H�4I�2��`���M�D(�m�j�!ݼ��C�66縂�m��؈&��}4e�!�F���;��B��"m%:���~���(p�
t3�f=�J���X��B�G��ɥ y�#M#Z�f�ЯD`���?�-�0�W�ף�������^�x��L7UD��F����P�]W�����RL��(��\6�뽵>`t༈D��G����!�HPQ�ڍ-*��gt��^�]e��M�� ��N%%�~>W��	Jqt��Y�,`��C��d��>;?g8�����ܘ��w�e����Ё}g`��]B��~hVe'[4���nZ;�o!սݰ��6��47^%��Y����>�c0���Yl���5���ϓjg0��`�=�́���lB��� ���t��4f�ʞ���*�-�x x}��4c F�o�X9�7�+ۍ2)���%�cG�t-���u���(�V2x_���U����ѧ�����8ce��9:�6]��>�(�	V�(z6Wgq�S�vd'���q���bm�5�)n+���j�G���6�b���9�yS���nS�^��e�jEb�OGk���:A����VX{c����wa)/�z4һ�G_��_A��30pX��578�8��O�� �63��'�AR.l�u��Gk������B�b=���&D3r���?����ُ.d��5�������S�XwA�ˡd�Ƃ�� �%�Thx��c�#�������pK%w��	��Q��$�21�[�q�п)�$>"�HW3� �7�qjP`F��\|>o��>��<��v��UV�ا�<Be��B��hJ����������9���卥��R)��-�d��Ԫ#��lt���#,�
�g8e(X ��p%�,�Ѳj��W�#��uɃ`y�|�누�"� �m�AhW���i6�ϐ#`�ap%���cb~�\M@g@按Di������'�vY4sp��[q�+1���Q��e4�{7#Uu�Գ�i��ZSx�6�;����V�\�����B<a�����Ƴ�����KK&a.�t�6��O��a!>-T��+���Fݓ��a'is	�"�ĬJ�p�����<��rr�ʓԀ7�o�g7"*��B��������8�j[:��*.W��XJ���B���P#�j�:�
�@˥s���*�ÔF\_�n�_~��BޢN�R%6[�n*�CW�f'���2�J敖d��&$�l,���g�i�sz��a���B<�f�X��I?.����Z�RE떺
�Ì�ńm��v2�[�m���Z����\�1¸g��FP�����t@)����~����m�иX�:�kn�s��m���(`4�,�	�䶺P���aX�a.@�m��neg�]RÆ�i�����i4љ�h�e^�!�1�}�������w�:<.���A�Q	����#����qr=Id��7�;�L�R(#�q��H��Ab�q��/f����s�&��������qh����}�hE�9౤Yd.Ju������n�g�A�,�}�cOoރ���$t_�2��ri���۾䇯���m:|%;��K���78�<���*�y�~�h���^�d����7�Ҵ@ u���i^%�<>���`����*�TBZ�����=���P[J
\@y��D�
nQj�%�����9(�� ��uZ��D�5z�(��a��c3f��q1op���&�{�^�����Nv`3�f��n�0������d�����C��"����8��kZ�ʇ8��p4TCo\����o�3������k�"b�B`����E��^�H��a�Cm�i$�e,>�x�7,4�?���D[:�ޞ�m^&�Q+�!w�\"�������Җ�#��B��GbϞ85ݩ���c�7`W�p@S�����.H~�֦���)[l����}_W�� n���F���~k��i%������M3�>��(�rnC4�M�.-M§���U@û�nÝ|�U9B$f�dXD�H\ �V���yX�j�>HA0��%���&q'TA��3��`�����.ak�Ev4��k���rjW��i�^n�X���מ�j�T����<p�����!%��.#��w��[aJe�0 ��mX:{p�v!&d�Y�zſ�ir���

��h�/���Y`���%Ti|A�� !9��ƭ)���H��{5�WH3ѹC����L�%�e�M���:,[��aPG�Ae������/��H�s����Sv�32P�pNQ��5�̣�'�HoC����f
&���ikD�r��H�!�xk-U\�ٴ��w�۵3�z*��V�𾓼�੬T@�:��Q,��]f� ;��J�l����|X�nc��0$_=��s��)f�&V�u��[}n隬�@o�j��F�t�	�I=�Z<qK��+�rN�l�g{����l�C�&1���)`�X-�XZ?���R�?u�h`�/@�O��|!�5�io�٧�1M>�0�emɷ���јɮ�E��L3�}q��8�ig�`g��!?��rD�M��f}�2��ʂ�C���	�ρ�U�Ϙ>?By�adA�w�t�}vi6�� ��5�a�<S�l�=�6�;Y&pB��ۣAt����P̳��MA+:�8'���1w"����@��+@w�qS��u�Tk�s�C���MhB�:�E1����Qd@������c�:s�T��zJǓ������H�'�`��\����%�ɳ�w����ౣ���3n�z����5�W!)j��Z���hct����Bj=<M���-�k�2�@�~p*ρ,w\���w�r�B�<�]��L�h����G>͎8Ԛ�B��)�`�����F���ן����� W���3�_zn��䅯#Ue��3Ҙ��,f�)+����K<��f~����F����!H�S���L�D����M���ZdO0
ڈ>�ȠDif�xA�w�H������QY��a|�!�(d�ݏ�Sah�ů-eؿ�rg�gI�R[$��0�b�8�b���N��5r���6h�/U�����fZ !ኪd՜��t���9�8�7*~4nsJ&��.��.C�z�l�-�`�H�B["&\����JPф���d߁众�����к��]���Ӽو:�4:�]'�D�5��D#M���&r\HM���KD:���!�x%�<$�.K��N�I �|	�-
����H���{e��c��
T�^{� 4k���E)�ѫ{A��,Ϛ����xV�6�Y��?7hB�O��K�L:?��Y�G�a��BObu�e�]8$���-������!�i������grn�M�r�\�W��l�	#G^�ퟞ_����S(���m��Yѷ��6�;􈓚���	kb��v����C����%bk��G�B���Ť��ash��C���?��B���[-��r�̦qT�+��j������`7̥e�u��j`�f/�m_�IR8]��}���|������I >�'9�iw�Y���������ۋ�	!S�B�z�wې�s�p}g�4�clV=��[a��_@�qG�������W�l�WOM��AߠG�!�@*I��uB�W!Lb��
�~�P9�Nhdjz��ʛ8=��
���M)�%��/Ƈh~�C;0���D��Y�B�b^fr�^DC�Kn���Y� �2U��rE@���fA�X@,|zgh�Q�x��4�%�A��u�Y�D
�]�R�
���Y+��F�/�Lȇ��ۮ��@��D����K�]2�M.�4����츷m�L���X��z5?�n^�E�R�;U�����r3�o��Eg9\�xs���$;�uC�z:R[�\j��'�7Esz����Oa���u�Fe��KI�g�
`�^%���N����bWN�I�u<�&�h��_�U~���y�@d6U��*Z�K��L�G<p�eCc�	�h�
��Yj���P�$���F}�$���.%-m^٬��Q�b�b[+��6�����..ٜ���̒L4R���R\�x�߃ l�A���(ܺ�xc�F�0�D�f+`�hh��CN\V���Ң��秌�r�G���Ԅ��ϭ�u:�b��9��*Tn�uR6��f�6S�qn)ݯz�e�v�?kNk� ld@Yc�{bH#���( ��iK|J.e�7vNf�k
xBr���@l���f�|K�8�.j��	P�~P����cd�`/E9��.��v,,�eI�'��6{�ζ���g���
�\���Z	.�vz
aO|��h��� T5�.�а���S����"A����o��3?�>���YD��W��rREv��V8"<[k�/�=v� )��]�9�V߿c0tͷt���o��QeX�`�U^$Vkyu�z�3�?ʲ�B��J�#"FX�,��e""��3�{�������x�[(�bl�8_1�� ��#��� |��<;IK�I�Uٍ7��`��W���gb��CUs{�{w�-����g�7��0�f�;�:u�\�)i��\(k���Q�S�#Y[GE��3^2� d�c��R�jza�`ݫ(l�
����1�>ZU|�õ.���d����7n��@��(�w��:<�3�<��IB�N%��00X�$�C�;��N�i�jP90�����o��Ǵ�吟�տ��n&1�͠�q�j
�����	v�:auy�(�ӚJc��%���յD6�">w��?�블y8�C n�U��Tӊ4��D2C8pJX���`�/�ț7�8�o�w���j�a�%�T�J��%H*)�����J���m����$��T����&!�S�MPS�Bŋ5��3`G�_Mk �f	G�z�t������,�>�g��;�wBX��gˣ4
��i`c�EĊ��T��N
]�}W� ��2۱K�
+yU�o{Zj��2~J�-�����<d������iG�FX�M��X�_�d(��>�6�4���g���#M�uh&g|�Y�1O^.�aHE}����P�9��/1�������3b����,�!�̫��_D���oWRlwn3����t�@W�'�H����K
�g�\���[�K`'�˗�ƕ�{bx�D��D�)$%�&f������x��ڊ2�m7�T_�i�֔�X��j��3eפ���X��T[�h�;L@�����l]B��jB9�Z�:֓������COdQ�7�)G��r":)E޲s�jb���0�S�j�Vo�3�QG���0��R�x�� �4
h�/[���9����ⓐ���#����M�>�Ú��jXH�6ys�.��͚��� k�W���춣�^�ɯ�j.k��ؽ��î�y���iXK���T[��0��|��RU4�w�S�EQ�D�\�j٪�����@!mr�&}-�M�媭mW���԰��S�/��)�1���!9E5�����m+k�rYϿ>��@_������ĉa���Aˮ6T20gޒ�G滧��`�T 4�2��]�����O���kPɨ}�,N�,�3����=L�,��D:�)�Ӊ��d�E�qX���$~��M���͖ˋ��7�jx��-7s�k������/�H}[�M�J�(�0�/?�r}�>��ein7��j]2��ž��OwP0���t�?�)�������3-�h�Z"
���@��׹�0�"�\�*⪇4x���#� ~rb��R�#�I9��PL	�փ�ȿ����~����\�0���wb��,,;}�]{��P�CK!RD \�t8k:��^�;�C���!�J�5g��O9`|��v�&4���n�㖎��RH ���<��I`���'I�{��8�=�1��"'7�����$���у��D�x���+� a�,��b��o��8G�R�6�x}�z���]X�w��a���I�n٤�|PP�n#�f�d�Q��U�,5�JW)������t��H���@�AmV-#�[�`Q�̧-��ӄA�L���l\8H�嫬�>5O��,:�� �Sf��I���p����T�_���a�T��:t�ve�g�'*�a!�$�� �ɨ��v����=�����y�a�:��ȉ'q��ȩ�BJժio�����g3PB.C3��f�"�x|r�u1��a���R�=�N�;�*���k��G-��7oI�BQ��q͞��$V1&�?r��_Ϲ���.��e���6�ǿ�X��~�t
���ԥ�#�tA!!����I ����UN�c>$�0 Ete�s�����G��N%'�r�O;�=�=�6	�GX8���l�)���g ^��ޏ�Ol(��r�!�
�60�_�l��\=P�Wu{4��Sx�;�~4�?� ����X��ȸ�֭'NЕ��	W�Ҋq���Թ	�%�A����al3���Z�`|�o;��j��i`>�'_`^;K�ˏ��JW��,���Ǡ�"�H�>	����O#��f������L~�M�a!4����7�s�yK�*'N:�ī�],��#��Z
#�|��<����s�-��PhZ�P*��A=�V�i�Z�v_g�4��� �����tu�)8�5�p)�jj�N���kE?�ފ�����&�\y7�E"�N�#����OȚRuez�t��:�:[�o�utƉV�"�>���k��Y�,�r{y��p�]楠Zr2o+'�f.����$1a�W@ߋ��َ�;���ӄ[��v[�����q8ѕ-s�CQ�=,�x��>�,��-�Ip3�qz�����NIV��S����q���%����V��o��5��6��m
��0� ��}���y��⍳�������'ƽss$�v}��^���t�c����.W d Hz�S��xh�P�w)	�e?P�Xy�lڇ�r����\��1�i�
�e�E/v1w�n������E=,ǂJڣ�t�fJ�>�}��މh��(��7x70�D��$2 B@�R�XPM|rTN�����Q�U\}�){������� ӣ+,)��2X�9X�S��TCFW8~aV�4[�-N��[�� B�# �Đ��y�1�ٷ���ڣ�J-��2�*@�r>����7:�~��}i��'��8H��.f,bc���ɯqAEh���k�� h2�/�.�����t�&�3͍�	ރ7k�T&w
^=a�*���J�wn?ߙ�l%���G'���ь.f�d0�P��5��"oPZ	%
!T ���9�v��x{x��9����Y������� ���ISdӉ�7K>��<7頴���l`�ǵϕ���7�IC]"��{ J�O6�> �Js��nn�P��+�,��*��W�fJ���(r�l/3�Z���%�3�%�so
e
\�jW�\�!Ӣޜ`�<�*�5���W�g�avr�w��c=އ9�0��oS��u��kz@����A/�B?��	���h=D����������3�ͳP?����<�wҧ��
!>g�IG���B�w=~Ԍ��6��y)�"������o���.D=r�/4i�@A$�:�]��
<�@z/$͏G	�"�Ʒq�|H �Wz�N�F��@�<��..��� ��dc}��KpL=��9Z4UB�X*�#_M�d��]Ip�6����u$�@v|��Ǚ�$�jTM45q�z����@� ���cM5���1͛{FZk�Nk��4�\�o�,��E���0�f�A�I8K $���1S����9Xw�\ܩO�m�ob���'kB����Fu�oj.�;ن�E��JqN��m� D�#�6/ CC)�d�A�h� x!�>�ȧ]Cis}8��EB���$��QG�v����;��|q;%ў0xT6kgO�����[woL(���h��f�����i�PO\��KӋ<:*叮�5��ȉ��l+�A?�A�����PN(R�ot�;�V]]�9`��
-H�Շ�T聄v���{�֚PA���NC�6�� ������EJ:��C��sU�fjJZ�v?�"��نFFu���\&�Z��%��M���V0N������<~%#4�*�ݔ���o1c �����3��m��5l�x�΀0�*%�9t�\8{s�h]�v�	%@Z���_ɧZe��4��\�$;��lT�z��l�9iHLP�T�fvzhS#��$T�F3�#�̥$�Q,S������J�N�9�u�/'W�>C�"���lX�D�v�T AN���]�bu*����\��aN����;�j.��z8�Or+�Pd���:@�q,��>J����}��S8g�|������	-���I3����]�e��/F�
2�		�e��]����	�0I垉���&�KT�-��w��Z���{�~h�����q�u��#T!���5ؖ,�,9H}��̹��Z�g���6�\1-�!�92:l�o��v8B�����\���&P���!�r91@Y�x��@���������Ęx]�>�����#BҘ��;�g���C%p�c
�]��H��n����2�3��X�8]zc�]]�0,�������<#䃟�&�\�=�F�Px�!���;��n!	h�l�ۣ������OI�6�f�LE������J���`>����?3��JSEw��j��tŀ��$�S��¥�k{�*��AO����Lb#-Y����/�?+1R�'lH�M�i���ԞYo� =�Y4F��:!�j�/q�
DW��@��k`�OD��}�4n' �]���m�	��
��6�ǀ�j9zF�v�P� l��@U �B�Z���s��r��
]ԓ�t>/fk�pr�1�P��- ŢJ�DT?<:&����� J�+���'��2�ryY6�2�E�T��~u�]��V�CZ�G䌨1৥�B�
�
 �TJ�>����T���Idi�辏h`�G�y��ex�7��Ee�9�.L��6a!���R�6��<bI%@�_Eɯ67\W�/s�W/WN��š?,��̿���۔�I$ԋB�m�6r>��ۥc+㧟F���:�;�U|

x�Uq��z80�%S߻u�x��~��n�q�-�J>����#E��.Z�⊩�5n��A��ugnp6�t��8������j��=_O�ȧ*�v�7g�4�Pk��Şܔ�e��{X��H���:0�����c3��,M|�W����ht48�Rbӿ��@0�b:+$�I�cQ<��AJ4���f�R�¿rˆ)��*m7�*�;ޤ��
T�JjU(Ȣ:?>M6R�f
ݷ[a�,�F��,������6!�%}7�1&;��B��'�1�za��䂪�w6�X�ƶͅ��;D փu�+���/#��rKe���v#��4l��
� ^����c�6ˆZ7tB{�y`���|R	�yj���,��������1M�q��,Vk��٢�e������մ\ҙN2ؖbV�����:�(�/��袐�q/+҃��v
��r'
�ŕ����x��̹��Ρ���+N���-�A�~rs�K��X�����pХदHh4]��5�5B�R��N�� m����Y���Y�H�l��s�s&Ot�y+�Gx�W\� �u�T|�$V�������0�;�uq ���vy&�9fㄾq��k���q���K�7bʁ���%1t `t�Oz�������$��!nRu,$6��p�y�V`�*|�X�D|M�L�ZW{ǧ^S������\WH������ '�����p�4n�9�F�Ś7�A%���(��]`yk��Y�,��/���$�e�[�4GI�4ϲ�qsP��[�xM�u���:l�O#&�]|�E:����'����L2Ս�%�S{�E;��-4@Q�G����.ܟ6�a�T1"����Od'ٟx��hs�~������Z��x��I#wBI���F*��d ���kW�	�y�w�������IJ��j�� Y�[ߖ J�^c���E�9NЮ�:-mw�����=�.k��E�[�Pl�Kr\ (��T$�Z4��Q������%)G�my=] ��8�><H[gm�z76+���t��C�w�J�V�+��o_�wE��j��C�ԯ,9a��P,ӌ/z$��o�i��yv�1�7(���um�p��eO���*N�����)	�HTz�gnj��,�c�1Jj��������@C�	��9�u���-I��pA��t�c��҃%��	�X1������A��F��G�E�I���`D�����^�*@�(�^;mﲒB����	#����иBpJ�<7�+�}�X���;r/&�uL;�Y�r���#��42�0�����۲��ْAPQ����E"Q����Pp�0���6<�������E�mk<�=�T���o�&	|Q�0�tM
=0��1�m]�X����@i�W��{Kc*�:J����[���*������v�_�N��&�f�]��~mC`��e��l/%=��3�-��1��*����h*6JaJ\, 1��l�%�ƗS^J��̘γ>߄�ef�*W�T��N�#>�~�0Q�*^Q��(���v}R�/�*wj/�?@	P�C�=/,�{<�Q�����d�Kui�����c�ю|%k�����c��&J�d���U��j5D� ��J�)��#ywJc�w	����$��9`/B����E�o���*���f8G9��R8���iu�@�_�{�&�	d̊���&��d�"{�w�u�WA�p��ْ�������~��旜��p��4@>��%3?j�@����2 ` �F�É=n�����5	�+	4��x�,�5�D��������%Hx�@���;r���hR��Ј�G0�n�������#�'WL:�O�a������jv �IHr�]>�Fȃ(��� �AÍ�d��f6�9��<
��f|6�)�c���K�(&o�bKC�EW�n�ę�S/��f5T��RI�5u��K� �t��S�.�c'R����
8E��GC��Ϯ2o����zW���c��s78�o�j�)����EG�g9.r6 �C�o��2 �r%%�D_�Βb�-�O
2�ps��Ii���~c!'Lh3�����?ۦȎ�9��R����%��;H�\�
�����N�$)�2��6�'�>��)�Tv_-_mKa�mD�=���z�[T�n됢���,�c�y=X�Nl�}»�6�Hdݙ|�g/7 �n�oS�I������ޝ% ��	�a5Z��T����>��a���u����M�(=� �/�~�_B.���7L�?���k��>��J���~�h�sc��|4����PU�k���q��SFծ���L���˫���xe}�GrϮ�k�7����Cf�[���%�\լ%VNg5o�O����rr�1��(���Lc�emt�Q�G�{r;Q�A�(���)��I
�Qf��F�^�e$�Ym=8nܾ���:?aˈ�Muw v�/����8KZ8�o�U�ڧdq����R�����`Z:�%��ܫ�a����k2��㿫z� �K-�$�ʚ@Yp"��7��O|���r�{�OJF�~N7�w��Ȏ��K,[��� ���Eܶ�����M���O_6�QP��Ţ�"Nk/�	㯲�o�ׁ���O_Gi�6G]�6y�,��pU~ZJ�K�.��VDo����qj�q�!S�rq)����p����(!X��~T��q&��0��SP/�-G�U 3��v�ݿ��)Hb6�?ʛ��G���g?*�4�Z\��u�?ɝ�-ss�R��,z!��-@�W�E�J�2����(�,����� ��P���b1�X=�q�Q�TL�j5w�-�#{�����$o_Pě m���`����:�����0�����&�;T�;���6���
��CX��(؊�H����r.���7���AI���7��gwX��`|T7^��%��u���c�^c�">�b����n��ʸ�W�{h��9����"2�l���1���P�U�oߎͤ[�7�=�Z��	-�;�:c��f&z1-%*�#��{�K�YN��("��T.�w_�~T� //�%~�R*���	ӊ?:5��q�|d��H�)6�>:� ��N�O�H�^��P&!��qb�v�����C̅p���^X���J��W��W�l����+�����#IE_XsZ�8m�xPH��D���G���|a/�{�����*����n�(0�bR��*߸�A������
�tfY�s��l�1�$�ȱ1����gg@E���~ov4��x�ޖ#����eRC>bV%�(�~A/�g���څ�R���,�����>�JW�?�vM'/F����>4A�W�yM��`#�t1�QS1��P,"�O�$=�Mk��GW��N�Q�X�p�~���V
(a3�����y�"��&���D�\�b��Kn���C�����E�����M���9�Z�@���	��=A���{���IZ.a���K`��X\b��p�R�ܱ)g����:�B���XV4p:�{ØZ����f��$B��٨qݺ��0���mj����^�X	w���&�����a,��a�o��rgIR��[]�����v!s�5�T4F��B���A�֍�n��-�ս	Z��@��c⻶D�������4��c�o�����1D�k�*��%au��-@�6�`A���5�D����ȊI��J���Fv�c!:lKb�z�U�X*Uq�5zɚ�#�YX��|u����
���(C��É^/��0��f,���������b���Ls	:��K�@|������e���Z����p�38����	�9H�Oَ��K߇y�T-TE�t����|�*Z<H;����!�G6�Q���yZU����]�΁6x$�&if�r�Na�2m��_�;�G���Kr�{�l�V���Y��$��a&&.�퓫�C6�w\��Թ�X;\
ą��Ӥ���f���Z���)�e�h8j���ޟs�F`7qU�
=m����`�l	��k�1�?����M &��94���]C���2����?2�����3�CBl�P�, 8k[�	�mp��h��Ua��V�i���l�
V�r�"��b�Յ����n����AOY�A���6�C����0'	v.�j�ݮ����A�ը�{���+��20'n��C��l�Ÿ�����]O�d�\"�$Ib^�Y��m�+1aQLa�2�4P���
[�����6f�|�5�T�m_)���?���%���9�m��/�����V����䟈O&�k�.L���˂��l�j�^<귥L��-��%�T��4���0T��6��b"Ly�@���;��;���_AA�3���a�7�	��ʹB�c�:w�|��Մ� \ܡ[0�D���~ڬtڠn��.5�V�+G I�2�|�&�!�Iy�xV������K
�A�dݖ��#���a��0"򻁐�8%9nױfz\��0��2�̵tx��{�p`q��/n`fOɭ����maAhU�����'m��jF�~QW����Ēu���U�`�?�Wz	�|��2t��`wO��9tKCC��h8Ԋ�V�g�:���r�T�l�CL���DN������ �	����:f�HD�E2�$�����MgR�5BxjYR1-���p/1�(%�� \������?L?�;��)�`lz��N�V�^�Z2��M��T�#GYL�����in�.�X�F��7�#ȡVN �-K�A�$
�w���=�|˼v�ꇨ�n���>1U+�ۀ��>�4�[���\&��o�X�>)�T�`�fЉ��o�^D���u�wI���(�w��-<�ӵm�⑭q��1�ɤ�b%��@]ilo=mB�$�W����:OE�@Y��qx�=���^���b!郪+��H8���k&���_��g7;ɰң�7��$bW.e�2�o��\�8��RD(���0���������x~�Q��������i}�#��	M̭��K��Jظ��X5�f�u�M�U �=f��'�"p!R�"��ì;���r��Y��EI_!�D��py�'�2FQT.��&l[��C�+N%��z#��[�po�5�����O3J����x��"OW�����ۥ��_� �H���f���|��^��6�gl��w�]�@���$�U:�@���8#���� W|��D8���W��Z�6�\ �!yӂ��15�S����L�P�	�y{��񸀾�����Y��ef�,���) i�3 ��Oٺ�������4^���d�I5�ʫ�v"�,���i|�����$_>74�f{���v����i�X�!�f�_�#��e�L��(�!��3DH��n[>T�3���Ӆ���4�x�A{�n�%iB��m�$c�����'�P�A�x�����������t?��E����2�hH�Ƕ��^쓇o!��SEK���Pϛ�!�1����{A�J:�ś������V˿S�pO��ʇ_�8��q-W����ͫ���t��9���Q�|rw�:�����f��DL�e�pG����I0��+Zݧ�Շ�p��`�ru��n��G)��݊�x�4�6VJ���v�!�Q�X��`��DV$�z�m"�e� ���o�q��ѩ����'�~Y-�o�V�9�3Or���R���gbR�!�ҙw�1MH��>�d�#��)��H���}�d��m�\��	V���$�l�*�d$�#����\���j���z��W?�d����Q}tZS����������t̓��;�f�Y��t>׳���Q<.Y��00�c�#_E�v^�&gDH�w���?�/���]��|˵��S��w����rYjY�*�%�z$�a&��"k�̨�@Ge��F�����}@�o,oȵ�c�&~��x�S�s��&8j��6�no�����*Qd��M2����-���R?ecRW�+� s�,��$%.���A�U����^���@��Ӛ.p�����:�����~yUK(5@�NE�#��-$��l�5�э�]1&�A�!wqw��iؼ���r�ֈ$�Ş�nɓ���m�!��q�5M���\����������V@rh�g�����<J�C�<!�Ռ�&sbOU,��L)<�-�,����'�&+���+G_l[^R�~�Ƚr0~r~�����q˦�"�7 `c�H1��
$��g�,z��<`�c�]���(B~�A^h �@A��ۏ�P^n;{/O���l^`nB��M@�4nݩ�^��o�QM�����U�>��#ia�J�W�$�}���%��W���4�����e���*�aX�"�*�&�d\�l`���2|ׅ�gN����Tՠ��6U�aC���ϋP7UsZ�k3�\I=�/u�ևF�#���+�	'DGH|b@S��~�ء�*˷4�qy��,\��.o�a��	��ނ��V��H���j;��a�i����]%���n(TK}`D�y��3��A�pn嬨BA��(*��c��/�E�+<|b���^DMWQ��0�F�kk����s~D�5����9�m�����X�^6,D�\�ɏ�Mk���)�����¡A�w�G�CJ��7Z��u�֌�Lk�H�'A�PY�]|f3&u�~)�LH�0��l'�*����n�w�@������� o-�?��Y�LMiE�>[���,z����Q#X��&Tf�N��Kz1���w��گA
����_� �|aKs�����w�^�u�d��>�;�9r�6q�?�(S\a�����/%���w���c�}{Ł	���ƽ��I�7z���Z�s�^��&s�l��'�z��W3g�������)��y<.ʫ��&D�`�`�=UD�ǫ	}C>֌�0��d	��+F��R�{	'��%X��L�<W�6W]��������ޣ|=as��*%��,8��������l{��=]�-Y�C�7�+�.�'���-�t�����Φ^߼��E��;ka�~��s%����.��z�{�?bK�b�|ܑ������r'c��F�=�p� ��{�8Ss3��4I�n)*-�(�����"�nb���K�U+G�>���3R�4yB3�&�k� Q0�BfS$�������Pfi\N(��j�&��*K��3I�!V�\fu�[�M�>P �(/�`��"l�Læ	&O��6�����Nh��ϴ��L&�'n�Z���:	� Ջm3�䳐{&�鰟0rΫ��\\4�����yr��w��缜�?� �f�!_N�kZ�<^zqj^�:i�غ�/��[�'�I��V�c��-�y�_�Tk��ZIAڭ��v�������`'Mn���bm�����B��©=����c���u1ަ_;4�<��N?�S���l[��m�뜣an B1�Ɵ�;+�+.�8�7،6dA>���D�����n��֭$��gq�&<Oz[�vn���zN��}�29�N��x�b�=Ϫ2��~R�V�%����YvR�~Cب�Դ�N�o�O�q���H���K"X%{b�$���0�zGʎ$��9m#�IT[���{��������K�!��m��M_]gk��a�{_y�E��=o�C\џ��U�|�>33�j
��Qp0��]?C
����,�x/���"5d�[���z��	�AM��P����.}�?�jB�`?u��ٱ�M�v�?4;�U��s0=��%/3��}LG-�K.�V �@��-�\����ш���pM�Vavw�e5�U�OjBd�Vjr�� ����uK!�
��;�5Y�mb}��%a����+)T�ic��[�fWW�������T� G ����?A8����Mvz�%��"���HSiD/g�
���������Z�oO��n,�t�� ����q�'��.�-���x�B�ʬ��՗�GR���׷�m�V��	r�k�j_KuOJM6;8G�#�x}+\P����WZ���Avڨq�_: �u�� �j8w�����Kڶ���$�w�E�݁EX�����C�PqQ�g�v�3���o��{b���GPCx��{F�����İ1�G�,Pu���\�Ӌ�Yl����b1�7�#VJ��1~|O�e����N��i ��v²��/�6�m�0\�#�8ʲ�QV~U�෶�m�A�?8�j��.o}DF�|�H{�[�]�t+C�y@�臍�0���������ϱ�#�UB�����AG7��v��D�2�ۏ���_�Ӓ���q�{�z@�(�#�:�$��Z�NΉ��Ns�����1�&�kF�`jǚ�"o�{C��ȲE���A��uy�����z����cÌµo���~+���#I�.���\�e�%�F@��eM�i�B/������?)��i����ap�tcg����u���q�˓���;��cxz�#�!�X�q��RB
���3�#+�L�s�8c������6��Jmӗ�k��}N���vC3�h+��}�7�B1�S��k^�h���R��Ƚ\(�ÿY(�#�ړeg�E��G@�S�jI��Q~\ʚ�7M*��/N~���a$w�"����CP��"��
2�ĚL=p\�s�����!�����p���u m���5���5T�����f���d{���$�8�&��MH}���Ǡ��j����,��A$M�j�� Ga��kt�n���:��#"�SEUC�D�vHTX��?�e�`@�W�Qҷ;���s^�ҝ�l�A�����Q�1a�]f�h�2�����2Ͽ$��U�N_��4��G���h�}ƀ
�ru��J^�����MW2j_/|)�w��u����{�Щ�W=4���8B[���n5B��lB0IK��՟TŪя�`|��%@��3��e�	�sVĺ#�8�K%� 3C2�4H������ܶR�)�r����Y>�/���"�c"F��f^l�'�-�e�HQ��t���?�V�	�+���n�a�W���/KW_�WS�۰)4����xmF���}��/�1̇��?�r�MևD`��