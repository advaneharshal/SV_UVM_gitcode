module top();
  initial
  begin
     $display("Shree Ganesha");
  end
endmodule
